module top (
            pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, 
            po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744;
assign w0 = ~pi0880 & ~pi2019;
assign w1 = ~pi0001 & pi2032;
assign w2 = ~pi0885 & ~pi2032;
assign w3 = ~pi0879 & ~pi0884;
assign w4 = ~pi0886 & ~pi0887;
assign w5 = ~pi0888 & ~pi0889;
assign w6 = ~pi0903 & w5;
assign w7 = w3 & w4;
assign w8 = w2 & w7;
assign w9 = w6 & w8;
assign w10 = ~w1 & ~w9;
assign w11 = pi0002 & pi2032;
assign w12 = pi0889 & ~pi2032;
assign w13 = ~w11 & ~w12;
assign w14 = pi0003 & pi2032;
assign w15 = pi0903 & ~pi2032;
assign w16 = ~w14 & ~w15;
assign w17 = pi0004 & pi2032;
assign w18 = pi0884 & ~pi2032;
assign w19 = ~w17 & ~w18;
assign w20 = ~pi0005 & pi2032;
assign w21 = ~w2 & ~w20;
assign w22 = pi0006 & pi2032;
assign w23 = pi0007 & pi2032;
assign w24 = pi0886 & ~pi2032;
assign w25 = ~w23 & ~w24;
assign w26 = pi0008 & pi2032;
assign w27 = pi0887 & ~pi2032;
assign w28 = ~w26 & ~w27;
assign w29 = pi0009 & pi2032;
assign w30 = pi0879 & ~pi2032;
assign w31 = ~w29 & ~w30;
assign w32 = pi0010 & pi2032;
assign w33 = pi0888 & ~pi2032;
assign w34 = ~w32 & ~w33;
assign w35 = pi0011 & pi2032;
assign w36 = pi0012 & pi2032;
assign w37 = pi0013 & pi2032;
assign w38 = pi0014 & pi2032;
assign w39 = pi0015 & pi2032;
assign w40 = pi0016 & pi2032;
assign w41 = pi0017 & pi2032;
assign w42 = pi1144 & ~pi2032;
assign w43 = ~w41 & ~w42;
assign w44 = pi0018 & pi2032;
assign w45 = pi1012 & ~pi2032;
assign w46 = ~w44 & ~w45;
assign w47 = pi0019 & pi2032;
assign w48 = pi1143 & ~pi2032;
assign w49 = ~w47 & ~w48;
assign w50 = pi0020 & pi2032;
assign w51 = pi1142 & ~pi2032;
assign w52 = ~w50 & ~w51;
assign w53 = pi0021 & pi2032;
assign w54 = pi1141 & ~pi2032;
assign w55 = ~w53 & ~w54;
assign w56 = pi0022 & pi2032;
assign w57 = pi1771 & ~pi2032;
assign w58 = ~w56 & ~w57;
assign w59 = pi0023 & pi2032;
assign w60 = pi1140 & ~pi2032;
assign w61 = ~w59 & ~w60;
assign w62 = pi0024 & pi2032;
assign w63 = pi1139 & ~pi2032;
assign w64 = ~w62 & ~w63;
assign w65 = pi0025 & pi2032;
assign w66 = pi0026 & pi2032;
assign w67 = pi0027 & pi2032;
assign w68 = pi0028 & pi2032;
assign w69 = pi0029 & pi2032;
assign w70 = pi0030 & pi2032;
assign w71 = pi0031 & pi2032;
assign w72 = pi0032 & pi2032;
assign w73 = pi0033 & pi2032;
assign w74 = pi0034 & pi2032;
assign w75 = pi0035 & pi2032;
assign w76 = pi0036 & pi2032;
assign w77 = pi0037 & pi2032;
assign w78 = ~pi1217 & ~pi2032;
assign w79 = ~w77 & ~w78;
assign w80 = pi0038 & pi2032;
assign w81 = ~pi1129 & ~pi2032;
assign w82 = ~w80 & ~w81;
assign w83 = pi0039 & pi2032;
assign w84 = ~pi1216 & ~pi2032;
assign w85 = ~w83 & ~w84;
assign w86 = pi0040 & pi2032;
assign w87 = ~pi1215 & ~pi2032;
assign w88 = ~w86 & ~w87;
assign w89 = pi0041 & pi2032;
assign w90 = ~pi1214 & ~pi2032;
assign w91 = ~w89 & ~w90;
assign w92 = pi0042 & pi2032;
assign w93 = ~pi1213 & ~pi2032;
assign w94 = ~w92 & ~w93;
assign w95 = pi0043 & pi2032;
assign w96 = ~pi1126 & ~pi2032;
assign w97 = ~w95 & ~w96;
assign w98 = pi0044 & pi2032;
assign w99 = ~pi1223 & ~pi2032;
assign w100 = ~w98 & ~w99;
assign w101 = pi0045 & pi2032;
assign w102 = ~pi1756 & ~pi2032;
assign w103 = ~w101 & ~w102;
assign w104 = pi0046 & pi2032;
assign w105 = ~pi1222 & ~pi2032;
assign w106 = ~w104 & ~w105;
assign w107 = pi0047 & pi2032;
assign w108 = ~pi1221 & ~pi2032;
assign w109 = ~w107 & ~w108;
assign w110 = pi0048 & pi2032;
assign w111 = ~pi1220 & ~pi2032;
assign w112 = ~w110 & ~w111;
assign w113 = pi0049 & pi2032;
assign w114 = ~pi1125 & ~pi2032;
assign w115 = ~w113 & ~w114;
assign w116 = pi0050 & pi2032;
assign w117 = ~pi1219 & ~pi2032;
assign w118 = ~w116 & ~w117;
assign w119 = pi0051 & pi2032;
assign w120 = ~pi1218 & ~pi2032;
assign w121 = ~w119 & ~w120;
assign w122 = pi0052 & pi2032;
assign w123 = ~pi1212 & ~pi2032;
assign w124 = ~w122 & ~w123;
assign w125 = pi0053 & pi2032;
assign w126 = pi0054 & pi2032;
assign w127 = pi0055 & pi2032;
assign w128 = pi0056 & pi2032;
assign w129 = pi0057 & pi2032;
assign w130 = ~pi0305 & ~pi2032;
assign w131 = ~w129 & ~w130;
assign w132 = pi0058 & pi2032;
assign w133 = ~pi0303 & ~pi2032;
assign w134 = ~w132 & ~w133;
assign w135 = pi0059 & pi2032;
assign w136 = ~pi0302 & ~pi2032;
assign w137 = ~w135 & ~w136;
assign w138 = pi0060 & pi2032;
assign w139 = ~pi0301 & ~pi2032;
assign w140 = ~w138 & ~w139;
assign w141 = pi0061 & pi2032;
assign w142 = ~pi0300 & ~pi2032;
assign w143 = ~w141 & ~w142;
assign w144 = pi0062 & pi2032;
assign w145 = ~pi0299 & ~pi2032;
assign w146 = ~w144 & ~w145;
assign w147 = pi0063 & pi2032;
assign w148 = ~pi0298 & ~pi2032;
assign w149 = ~w147 & ~w148;
assign w150 = pi0064 & pi2032;
assign w151 = ~pi0308 & ~pi2032;
assign w152 = ~w150 & ~w151;
assign w153 = pi0065 & pi2032;
assign w154 = ~pi0297 & ~pi2032;
assign w155 = ~w153 & ~w154;
assign w156 = pi0066 & pi2032;
assign w157 = ~pi0296 & ~pi2032;
assign w158 = ~w156 & ~w157;
assign w159 = pi0067 & pi2032;
assign w160 = ~pi0321 & ~pi2032;
assign w161 = ~w159 & ~w160;
assign w162 = pi0068 & pi2032;
assign w163 = ~pi0317 & ~pi2032;
assign w164 = ~w162 & ~w163;
assign w165 = pi0069 & pi2032;
assign w166 = ~pi0315 & ~pi2032;
assign w167 = ~w165 & ~w166;
assign w168 = pi0070 & pi2032;
assign w169 = ~pi0313 & ~pi2032;
assign w170 = ~w168 & ~w169;
assign w171 = pi0071 & pi2032;
assign w172 = ~pi0319 & ~pi2032;
assign w173 = ~w171 & ~w172;
assign w174 = pi0072 & pi2032;
assign w175 = ~pi0311 & ~pi2032;
assign w176 = ~w174 & ~w175;
assign w177 = pi0073 & pi2032;
assign w178 = ~pi0245 & ~pi2032;
assign w179 = ~w177 & ~w178;
assign w180 = pi0074 & pi2032;
assign w181 = ~pi0244 & ~pi2032;
assign w182 = ~w180 & ~w181;
assign w183 = pi0075 & pi2032;
assign w184 = ~pi0258 & ~pi2032;
assign w185 = ~w183 & ~w184;
assign w186 = pi0076 & pi2032;
assign w187 = ~pi0256 & ~pi2032;
assign w188 = ~w186 & ~w187;
assign w189 = pi0077 & pi2032;
assign w190 = ~pi0421 & ~pi2032;
assign w191 = ~w189 & ~w190;
assign w192 = pi0078 & pi2032;
assign w193 = ~pi0419 & ~pi2032;
assign w194 = ~w192 & ~w193;
assign w195 = pi0079 & pi2032;
assign w196 = ~pi0422 & ~pi2032;
assign w197 = ~w195 & ~w196;
assign w198 = pi0080 & pi2032;
assign w199 = ~pi0417 & ~pi2032;
assign w200 = ~w198 & ~w199;
assign w201 = pi0081 & pi2032;
assign w202 = ~pi0416 & ~pi2032;
assign w203 = ~w201 & ~w202;
assign w204 = pi0082 & pi2032;
assign w205 = ~pi0415 & ~pi2032;
assign w206 = ~w204 & ~w205;
assign w207 = pi0083 & pi2032;
assign w208 = ~pi0414 & ~pi2032;
assign w209 = ~w207 & ~w208;
assign w210 = pi0084 & pi2032;
assign w211 = ~pi0420 & ~pi2032;
assign w212 = ~w210 & ~w211;
assign w213 = pi0085 & pi2032;
assign w214 = ~pi0418 & ~pi2032;
assign w215 = ~w213 & ~w214;
assign w216 = pi0086 & pi2032;
assign w217 = ~pi0413 & ~pi2032;
assign w218 = ~w216 & ~w217;
assign w219 = pi0087 & pi2032;
assign w220 = ~pi0427 & ~pi2032;
assign w221 = ~w219 & ~w220;
assign w222 = pi0088 & pi2032;
assign w223 = ~pi0426 & ~pi2032;
assign w224 = ~w222 & ~w223;
assign w225 = pi0089 & pi2032;
assign w226 = ~pi0425 & ~pi2032;
assign w227 = ~w225 & ~w226;
assign w228 = pi0090 & pi2032;
assign w229 = ~pi0424 & ~pi2032;
assign w230 = ~w228 & ~w229;
assign w231 = pi0091 & pi2032;
assign w232 = ~pi0423 & ~pi2032;
assign w233 = ~w231 & ~w232;
assign w234 = pi0092 & pi2032;
assign w235 = ~pi0345 & ~pi2032;
assign w236 = ~w234 & ~w235;
assign w237 = pi0093 & pi2032;
assign w238 = ~pi0337 & ~pi2032;
assign w239 = ~w237 & ~w238;
assign w240 = pi0094 & pi2032;
assign w241 = ~pi0340 & ~pi2032;
assign w242 = ~w240 & ~w241;
assign w243 = pi0095 & pi2032;
assign w244 = ~pi0351 & ~pi2032;
assign w245 = ~w243 & ~w244;
assign w246 = pi0096 & pi2032;
assign w247 = ~pi0352 & ~pi2032;
assign w248 = ~w246 & ~w247;
assign w249 = pi0097 & pi2032;
assign w250 = pi0098 & pi2032;
assign w251 = pi0099 & pi2032;
assign w252 = pi0100 & pi2032;
assign w253 = pi0101 & pi2032;
assign w254 = pi0102 & pi2032;
assign w255 = pi0103 & pi2032;
assign w256 = pi0104 & pi2032;
assign w257 = pi0105 & pi2032;
assign w258 = pi0106 & pi2032;
assign w259 = pi0107 & pi2032;
assign w260 = pi0108 & pi2032;
assign w261 = pi0109 & pi2032;
assign w262 = pi0110 & pi2032;
assign w263 = pi0111 & pi2032;
assign w264 = pi0112 & pi2032;
assign w265 = pi0113 & pi2032;
assign w266 = pi0114 & pi2032;
assign w267 = pi0115 & pi2032;
assign w268 = pi0116 & pi2032;
assign w269 = pi0117 & pi2032;
assign w270 = ~pi0435 & ~pi2032;
assign w271 = ~w269 & ~w270;
assign w272 = pi0118 & pi2032;
assign w273 = ~pi0434 & ~pi2032;
assign w274 = ~w272 & ~w273;
assign w275 = pi0119 & pi2032;
assign w276 = ~pi0455 & ~pi2032;
assign w277 = ~w275 & ~w276;
assign w278 = pi0120 & pi2032;
assign w279 = ~pi0433 & ~pi2032;
assign w280 = ~w278 & ~w279;
assign w281 = pi0121 & pi2032;
assign w282 = ~pi0432 & ~pi2032;
assign w283 = ~w281 & ~w282;
assign w284 = pi0122 & pi2032;
assign w285 = ~pi0431 & ~pi2032;
assign w286 = ~w284 & ~w285;
assign w287 = pi0123 & pi2032;
assign w288 = ~pi0457 & ~pi2032;
assign w289 = ~w287 & ~w288;
assign w290 = pi0124 & pi2032;
assign w291 = ~pi0430 & ~pi2032;
assign w292 = ~w290 & ~w291;
assign w293 = pi0125 & pi2032;
assign w294 = ~pi0429 & ~pi2032;
assign w295 = ~w293 & ~w294;
assign w296 = pi0126 & pi2032;
assign w297 = ~pi0428 & ~pi2032;
assign w298 = ~w296 & ~w297;
assign w299 = pi0127 & pi2032;
assign w300 = ~pi0440 & ~pi2032;
assign w301 = ~w299 & ~w300;
assign w302 = pi0128 & pi2032;
assign w303 = ~pi0439 & ~pi2032;
assign w304 = ~w302 & ~w303;
assign w305 = pi0129 & pi2032;
assign w306 = ~pi0454 & ~pi2032;
assign w307 = ~w305 & ~w306;
assign w308 = pi0130 & pi2032;
assign w309 = ~pi0438 & ~pi2032;
assign w310 = ~w308 & ~w309;
assign w311 = pi0131 & pi2032;
assign w312 = ~pi0437 & ~pi2032;
assign w313 = ~w311 & ~w312;
assign w314 = pi0132 & pi2032;
assign w315 = ~pi0436 & ~pi2032;
assign w316 = ~w314 & ~w315;
assign w317 = pi0133 & pi2032;
assign w318 = ~pi0338 & ~pi2032;
assign w319 = ~w317 & ~w318;
assign w320 = pi0134 & pi2032;
assign w321 = ~pi0339 & ~pi2032;
assign w322 = ~w320 & ~w321;
assign w323 = pi0135 & pi2032;
assign w324 = ~pi0350 & ~pi2032;
assign w325 = ~w323 & ~w324;
assign w326 = pi0136 & pi2032;
assign w327 = ~pi0349 & ~pi2032;
assign w328 = ~w326 & ~w327;
assign w329 = pi0137 & pi2032;
assign w330 = ~pi0271 & ~pi2032;
assign w331 = ~w329 & ~w330;
assign w332 = pi0138 & pi2032;
assign w333 = ~pi0270 & ~pi2032;
assign w334 = ~w332 & ~w333;
assign w335 = pi0139 & pi2032;
assign w336 = ~pi0273 & ~pi2032;
assign w337 = ~w335 & ~w336;
assign w338 = pi0140 & pi2032;
assign w339 = ~pi0272 & ~pi2032;
assign w340 = ~w338 & ~w339;
assign w341 = pi0141 & pi2032;
assign w342 = ~pi0267 & ~pi2032;
assign w343 = ~w341 & ~w342;
assign w344 = pi0142 & pi2032;
assign w345 = ~pi0266 & ~pi2032;
assign w346 = ~w344 & ~w345;
assign w347 = pi0143 & pi2032;
assign w348 = ~pi0265 & ~pi2032;
assign w349 = ~w347 & ~w348;
assign w350 = pi0144 & pi2032;
assign w351 = ~pi0264 & ~pi2032;
assign w352 = ~w350 & ~w351;
assign w353 = pi0145 & pi2032;
assign w354 = ~pi0269 & ~pi2032;
assign w355 = ~w353 & ~w354;
assign w356 = pi0146 & pi2032;
assign w357 = ~pi0268 & ~pi2032;
assign w358 = ~w356 & ~w357;
assign w359 = pi0147 & pi2032;
assign w360 = ~pi0279 & ~pi2032;
assign w361 = ~w359 & ~w360;
assign w362 = pi0148 & pi2032;
assign w363 = ~pi0278 & ~pi2032;
assign w364 = ~w362 & ~w363;
assign w365 = pi0149 & pi2032;
assign w366 = ~pi0277 & ~pi2032;
assign w367 = ~w365 & ~w366;
assign w368 = pi0150 & pi2032;
assign w369 = ~pi0276 & ~pi2032;
assign w370 = ~w368 & ~w369;
assign w371 = pi0151 & pi2032;
assign w372 = ~pi0275 & ~pi2032;
assign w373 = ~w371 & ~w372;
assign w374 = pi0152 & pi2032;
assign w375 = ~pi0274 & ~pi2032;
assign w376 = ~w374 & ~w375;
assign w377 = pi0153 & pi2032;
assign w378 = ~pi0241 & ~pi2032;
assign w379 = ~w377 & ~w378;
assign w380 = pi0154 & pi2032;
assign w381 = ~pi0240 & ~pi2032;
assign w382 = ~w380 & ~w381;
assign w383 = pi0155 & pi2032;
assign w384 = ~pi0253 & ~pi2032;
assign w385 = ~w383 & ~w384;
assign w386 = pi0156 & pi2032;
assign w387 = ~pi0252 & ~pi2032;
assign w388 = ~w386 & ~w387;
assign w389 = pi0157 & pi2032;
assign w390 = ~pi0287 & ~pi2032;
assign w391 = ~w389 & ~w390;
assign w392 = pi0158 & pi2032;
assign w393 = ~pi0289 & ~pi2032;
assign w394 = ~w392 & ~w393;
assign w395 = pi0159 & pi2032;
assign w396 = ~pi0285 & ~pi2032;
assign w397 = ~w395 & ~w396;
assign w398 = pi0160 & pi2032;
assign w399 = ~pi0288 & ~pi2032;
assign w400 = ~w398 & ~w399;
assign w401 = pi0161 & pi2032;
assign w402 = ~pi0286 & ~pi2032;
assign w403 = ~w401 & ~w402;
assign w404 = pi0162 & pi2032;
assign w405 = ~pi0284 & ~pi2032;
assign w406 = ~w404 & ~w405;
assign w407 = pi0163 & pi2032;
assign w408 = ~pi0283 & ~pi2032;
assign w409 = ~w407 & ~w408;
assign w410 = pi0164 & pi2032;
assign w411 = ~pi0282 & ~pi2032;
assign w412 = ~w410 & ~w411;
assign w413 = pi0165 & pi2032;
assign w414 = ~pi0281 & ~pi2032;
assign w415 = ~w413 & ~w414;
assign w416 = pi0166 & pi2032;
assign w417 = ~pi0280 & ~pi2032;
assign w418 = ~w416 & ~w417;
assign w419 = pi0167 & pi2032;
assign w420 = ~pi0295 & ~pi2032;
assign w421 = ~w419 & ~w420;
assign w422 = pi0168 & pi2032;
assign w423 = ~pi0294 & ~pi2032;
assign w424 = ~w422 & ~w423;
assign w425 = pi0169 & pi2032;
assign w426 = ~pi0293 & ~pi2032;
assign w427 = ~w425 & ~w426;
assign w428 = pi0170 & pi2032;
assign w429 = ~pi0292 & ~pi2032;
assign w430 = ~w428 & ~w429;
assign w431 = pi0171 & pi2032;
assign w432 = ~pi0291 & ~pi2032;
assign w433 = ~w431 & ~w432;
assign w434 = pi0172 & pi2032;
assign w435 = ~pi0290 & ~pi2032;
assign w436 = ~w434 & ~w435;
assign w437 = pi0173 & pi2032;
assign w438 = ~pi0243 & ~pi2032;
assign w439 = ~w437 & ~w438;
assign w440 = pi0174 & pi2032;
assign w441 = ~pi0242 & ~pi2032;
assign w442 = ~w440 & ~w441;
assign w443 = pi0175 & pi2032;
assign w444 = ~pi0255 & ~pi2032;
assign w445 = ~w443 & ~w444;
assign w446 = pi0176 & pi2032;
assign w447 = ~pi0254 & ~pi2032;
assign w448 = ~w446 & ~w447;
assign w449 = pi0177 & pi2032;
assign w450 = ~pi0320 & ~pi2032;
assign w451 = ~w449 & ~w450;
assign w452 = pi0178 & pi2032;
assign w453 = ~pi0316 & ~pi2032;
assign w454 = ~w452 & ~w453;
assign w455 = pi0179 & pi2032;
assign w456 = ~pi0314 & ~pi2032;
assign w457 = ~w455 & ~w456;
assign w458 = pi0180 & pi2032;
assign w459 = ~pi0312 & ~pi2032;
assign w460 = ~w458 & ~w459;
assign w461 = pi0181 & pi2032;
assign w462 = ~pi0318 & ~pi2032;
assign w463 = ~w461 & ~w462;
assign w464 = pi0182 & pi2032;
assign w465 = ~pi0310 & ~pi2032;
assign w466 = ~w464 & ~w465;
assign w467 = pi0183 & pi2032;
assign w468 = ~pi0309 & ~pi2032;
assign w469 = ~w467 & ~w468;
assign w470 = pi0184 & pi2032;
assign w471 = ~pi0307 & ~pi2032;
assign w472 = ~w470 & ~w471;
assign w473 = pi0185 & pi2032;
assign w474 = ~pi0306 & ~pi2032;
assign w475 = ~w473 & ~w474;
assign w476 = pi0186 & pi2032;
assign w477 = ~pi0304 & ~pi2032;
assign w478 = ~w476 & ~w477;
assign w479 = pi0187 & pi2032;
assign w480 = ~pi0327 & ~pi2032;
assign w481 = ~w479 & ~w480;
assign w482 = pi0188 & pi2032;
assign w483 = ~pi0326 & ~pi2032;
assign w484 = ~w482 & ~w483;
assign w485 = pi0189 & pi2032;
assign w486 = ~pi0325 & ~pi2032;
assign w487 = ~w485 & ~w486;
assign w488 = pi0200 & pi2032;
assign w489 = ~pi0324 & ~pi2032;
assign w490 = ~w488 & ~w489;
assign w491 = pi0190 & pi2056;
assign w492 = pi0209 & ~pi2056;
assign w493 = ~w491 & ~w492;
assign w494 = pi0191 & pi2059;
assign w495 = pi0209 & ~pi2059;
assign w496 = ~w494 & ~w495;
assign w497 = pi0192 & pi2057;
assign w498 = pi0209 & ~pi2057;
assign w499 = ~w497 & ~w498;
assign w500 = pi0193 & pi2058;
assign w501 = pi0209 & ~pi2058;
assign w502 = ~w500 & ~w501;
assign w503 = pi0194 & pi2056;
assign w504 = pi0228 & ~pi2056;
assign w505 = ~w503 & ~w504;
assign w506 = pi0195 & pi2059;
assign w507 = pi0228 & ~pi2059;
assign w508 = ~w506 & ~w507;
assign w509 = pi0196 & pi2057;
assign w510 = pi0228 & ~pi2057;
assign w511 = ~w509 & ~w510;
assign w512 = pi0197 & pi2058;
assign w513 = pi0228 & ~pi2058;
assign w514 = ~w512 & ~w513;
assign w515 = ~pi1167 & ~pi1987;
assign w516 = pi1167 & pi1987;
assign w517 = ~pi1166 & ~pi2140;
assign w518 = ~w516 & w517;
assign w519 = pi1903 & ~w515;
assign w520 = ~w518 & w519;
assign w521 = pi1035 & ~w520;
assign w522 = ~w520 & w9594;
assign w523 = (~pi0198 & w520) | (~pi0198 & w9596) | (w520 & w9596);
assign w524 = ~pi2247 & ~w523;
assign w525 = ~pi1180 & ~pi2005;
assign w526 = pi1180 & pi2005;
assign w527 = ~pi1179 & ~pi2138;
assign w528 = ~w526 & w527;
assign w529 = pi1904 & ~w525;
assign w530 = ~w528 & w529;
assign w531 = pi1176 & ~w530;
assign w532 = ~w530 & w9597;
assign w533 = (~pi0199 & w530) | (~pi0199 & w9599) | (w530 & w9599);
assign w534 = ~pi2249 & ~w533;
assign w535 = pi0328 & pi2032;
assign w536 = ~pi0323 & ~pi2032;
assign w537 = ~w535 & ~w536;
assign w538 = ~pi1184 & ~pi2004;
assign w539 = pi1184 & pi2004;
assign w540 = ~pi1131 & ~pi2139;
assign w541 = ~w539 & w540;
assign w542 = pi1907 & ~w538;
assign w543 = ~w541 & w542;
assign w544 = pi1164 & ~w543;
assign w545 = ~w543 & w9600;
assign w546 = (~pi0201 & w543) | (~pi0201 & w9602) | (w543 & w9602);
assign w547 = ~pi2246 & ~w546;
assign w548 = ~pi1174 & ~pi1988;
assign w549 = pi1174 & pi1988;
assign w550 = ~pi1173 & ~pi2158;
assign w551 = ~w549 & w550;
assign w552 = pi1908 & ~w548;
assign w553 = ~w551 & w552;
assign w554 = pi1169 & ~w553;
assign w555 = ~w553 & w9603;
assign w556 = (~pi0202 & w553) | (~pi0202 & w9605) | (w553 & w9605);
assign w557 = ~pi2248 & ~w556;
assign w558 = ~pi1847 & ~pi2006;
assign w559 = pi1847 & pi2006;
assign w560 = ~pi1873 & ~pi2141;
assign w561 = ~w559 & w560;
assign w562 = pi1909 & ~w558;
assign w563 = ~w561 & w562;
assign w564 = pi1839 & ~w563;
assign w565 = ~w563 & w9606;
assign w566 = (~pi0203 & w563) | (~pi0203 & w9608) | (w563 & w9608);
assign w567 = ~pi2250 & ~w566;
assign w568 = ~pi1842 & ~pi2007;
assign w569 = pi1842 & pi2007;
assign w570 = ~pi1841 & ~pi2159;
assign w571 = ~w569 & w570;
assign w572 = pi1910 & ~w568;
assign w573 = ~w571 & w572;
assign w574 = pi1838 & ~w573;
assign w575 = ~w573 & w9609;
assign w576 = (~pi0204 & w573) | (~pi0204 & w9611) | (w573 & w9611);
assign w577 = ~pi2251 & ~w576;
assign w578 = pi0205 & pi2056;
assign w579 = pi0331 & ~pi2056;
assign w580 = ~w578 & ~w579;
assign w581 = pi0206 & pi2059;
assign w582 = pi0331 & ~pi2059;
assign w583 = ~w581 & ~w582;
assign w584 = pi0207 & pi2057;
assign w585 = pi0331 & ~pi2057;
assign w586 = ~w584 & ~w585;
assign w587 = pi0208 & pi2058;
assign w588 = pi0331 & ~pi2058;
assign w589 = ~w587 & ~w588;
assign w590 = pi0210 & pi2056;
assign w591 = pi0456 & ~pi2056;
assign w592 = ~w590 & ~w591;
assign w593 = pi0211 & pi2059;
assign w594 = pi0456 & ~pi2059;
assign w595 = ~w593 & ~w594;
assign w596 = pi0212 & pi2057;
assign w597 = pi0456 & ~pi2057;
assign w598 = ~w596 & ~w597;
assign w599 = pi0213 & pi2058;
assign w600 = pi0456 & ~pi2058;
assign w601 = ~w599 & ~w600;
assign w602 = pi0885 & pi1930;
assign w603 = ~pi1076 & w602;
assign w604 = ~pi1020 & ~pi1165;
assign w605 = ~pi0353 & w604;
assign w606 = w603 & ~w605;
assign w607 = w606 & w2282;
assign w608 = (w606 & w9612) | (w606 & w9613) | (w9612 & w9613);
assign w609 = ~w607 & w608;
assign w610 = ~pi0215 & pi0238;
assign w611 = ~pi1171 & ~pi1789;
assign w612 = ~pi0354 & w611;
assign w613 = pi0886 & pi1930;
assign w614 = ~pi1077 & w613;
assign w615 = ~w612 & w614;
assign w616 = w615 & w9614;
assign w617 = (pi1169 & ~w615) | (pi1169 & w9615) | (~w615 & w9615);
assign w618 = ~w616 & ~w617;
assign w619 = (~pi0215 & ~w615) | (~pi0215 & w9616) | (~w615 & w9616);
assign w620 = ~w618 & ~w619;
assign w621 = pi0888 & pi1930;
assign w622 = ~pi1080 & w621;
assign w623 = ~pi1832 & ~pi1840;
assign w624 = ~pi0260 & w623;
assign w625 = w622 & ~w624;
assign w626 = w625 & w863;
assign w627 = (w625 & w9617) | (w625 & w9618) | (w9617 & w9618);
assign w628 = ~w626 & w627;
assign w629 = pi0884 & pi1930;
assign w630 = ~pi1075 & w629;
assign w631 = ~pi1130 & ~pi1183;
assign w632 = ~pi0261 & w631;
assign w633 = w630 & ~w632;
assign w634 = w633 & w813;
assign w635 = (w633 & w9619) | (w633 & w9620) | (w9619 & w9620);
assign w636 = ~w634 & w635;
assign w637 = pi0887 & pi1930;
assign w638 = ~pi1078 & w637;
assign w639 = ~pi1178 & ~pi1777;
assign w640 = ~pi0262 & w639;
assign w641 = w638 & ~w640;
assign w642 = w641 & w725;
assign w643 = (w641 & w9621) | (w641 & w9622) | (w9621 & w9622);
assign w644 = ~w642 & w643;
assign w645 = pi0879 & pi1930;
assign w646 = ~pi1079 & w645;
assign w647 = ~pi1845 & ~pi1846;
assign w648 = ~pi0263 & w647;
assign w649 = w646 & ~w648;
assign w650 = w649 & w773;
assign w651 = (w649 & w9623) | (w649 & w9624) | (w9623 & w9624);
assign w652 = ~w650 & w651;
assign w653 = w625 & w9626;
assign w654 = (w625 & w9627) | (w625 & w9628) | (w9627 & w9628);
assign w655 = ~w653 & w654;
assign w656 = w633 & w9630;
assign w657 = (w633 & w9631) | (w633 & w9632) | (w9631 & w9632);
assign w658 = ~w656 & w657;
assign w659 = w641 & w9634;
assign w660 = (w641 & w9635) | (w641 & w9636) | (w9635 & w9636);
assign w661 = ~w659 & w660;
assign w662 = w649 & w9638;
assign w663 = (w649 & w9639) | (w649 & w9640) | (w9639 & w9640);
assign w664 = ~w662 & w663;
assign w665 = ~pi0224 & ~w625;
assign w666 = (pi1838 & ~w625) | (pi1838 & w9641) | (~w625 & w9641);
assign w667 = ~w665 & w666;
assign w668 = ~pi0225 & ~w633;
assign w669 = (pi1164 & ~w633) | (pi1164 & w9642) | (~w633 & w9642);
assign w670 = ~w668 & w669;
assign w671 = ~pi0226 & ~w649;
assign w672 = (pi1839 & ~w649) | (pi1839 & w9643) | (~w649 & w9643);
assign w673 = ~w671 & w672;
assign w674 = ~pi0227 & ~w641;
assign w675 = (pi1176 & ~w641) | (pi1176 & w9644) | (~w641 & w9644);
assign w676 = ~w674 & w675;
assign w677 = ~pi0229 & ~pi0838;
assign w678 = ~pi2238 & pi2239;
assign w679 = pi2240 & w678;
assign w680 = ~pi2241 & ~pi2242;
assign w681 = pi2202 & pi2203;
assign w682 = ~pi2131 & ~pi2201;
assign w683 = w681 & w682;
assign w684 = pi2132 & w683;
assign w685 = w679 & w680;
assign w686 = w684 & w685;
assign w687 = ~w677 & ~w686;
assign w688 = ~pi0230 & ~pi0839;
assign w689 = ~w686 & ~w688;
assign w690 = pi0231 & pi2059;
assign w691 = pi0640 & ~pi2059;
assign w692 = ~w690 & ~w691;
assign w693 = pi0640 & pi2060;
assign w694 = pi0232 & ~pi2060;
assign w695 = ~w693 & ~w694;
assign w696 = pi0233 & pi2058;
assign w697 = pi0640 & ~pi2058;
assign w698 = ~w696 & ~w697;
assign w699 = pi0234 & pi2056;
assign w700 = pi0640 & ~pi2056;
assign w701 = ~w699 & ~w700;
assign w702 = pi0235 & pi2057;
assign w703 = pi0640 & ~pi2057;
assign w704 = ~w702 & ~w703;
assign w705 = ~pi0236 & ~w606;
assign w706 = (pi1035 & ~w606) | (pi1035 & w9645) | (~w606 & w9645);
assign w707 = ~w705 & w706;
assign w708 = w606 & w9647;
assign w709 = (w606 & w9648) | (w606 & w9649) | (w9648 & w9649);
assign w710 = ~w708 & w709;
assign w711 = ~pi0238 & ~w615;
assign w712 = w617 & ~w711;
assign w713 = pi0239 & ~w618;
assign w714 = pi0215 & pi0238;
assign w715 = ~pi0239 & w714;
assign w716 = w615 & w9650;
assign w717 = ~w713 & ~w716;
assign w718 = w637 & w9651;
assign w719 = ~pi1178 & pi1777;
assign w720 = w718 & w719;
assign w721 = ~pi0218 & ~pi0227;
assign w722 = pi1758 & w721;
assign w723 = ~pi0218 & pi0227;
assign w724 = pi1461 & w723;
assign w725 = pi0218 & pi0227;
assign w726 = pi1510 & w725;
assign w727 = pi0218 & ~pi0227;
assign w728 = pi1486 & w727;
assign w729 = ~w722 & ~w724;
assign w730 = ~w726 & ~w728;
assign w731 = w729 & w730;
assign w732 = (pi1176 & ~w637) | (pi1176 & w9652) | (~w637 & w9652);
assign w733 = ~pi0240 & w732;
assign w734 = pi1178 & ~pi1777;
assign w735 = w718 & w734;
assign w736 = pi1795 & w723;
assign w737 = pi1775 & w727;
assign w738 = pi1709 & w721;
assign w739 = pi1761 & w725;
assign w740 = ~w736 & ~w737;
assign w741 = ~w738 & ~w739;
assign w742 = w740 & w741;
assign w743 = w735 & ~w742;
assign w744 = (~w733 & w731) | (~w733 & w9653) | (w731 & w9653);
assign w745 = ~w743 & w744;
assign w746 = pi1704 & w721;
assign w747 = pi1518 & w725;
assign w748 = pi1494 & w727;
assign w749 = pi1470 & w723;
assign w750 = ~w746 & ~w747;
assign w751 = ~w748 & ~w749;
assign w752 = w750 & w751;
assign w753 = ~pi0241 & w732;
assign w754 = pi1711 & w721;
assign w755 = pi1529 & w725;
assign w756 = pi1481 & w723;
assign w757 = pi1505 & w727;
assign w758 = ~w754 & ~w755;
assign w759 = ~w756 & ~w757;
assign w760 = w758 & w759;
assign w761 = w735 & ~w760;
assign w762 = (~w753 & w752) | (~w753 & w9654) | (w752 & w9654);
assign w763 = ~w761 & w762;
assign w764 = w645 & w9655;
assign w765 = pi1845 & ~pi1846;
assign w766 = w764 & w765;
assign w767 = pi0219 & ~pi0226;
assign w768 = pi1560 & w767;
assign w769 = ~pi0219 & pi0226;
assign w770 = pi1535 & w769;
assign w771 = ~pi0219 & ~pi0226;
assign w772 = pi1102 & w771;
assign w773 = pi0219 & pi0226;
assign w774 = pi1584 & w773;
assign w775 = ~w768 & ~w770;
assign w776 = ~w772 & ~w774;
assign w777 = w775 & w776;
assign w778 = (pi1839 & ~w645) | (pi1839 & w9656) | (~w645 & w9656);
assign w779 = ~pi0242 & w778;
assign w780 = ~pi1845 & pi1846;
assign w781 = w764 & w780;
assign w782 = pi1552 & w769;
assign w783 = pi1576 & w767;
assign w784 = pi1601 & w773;
assign w785 = pi1724 & w771;
assign w786 = ~w782 & ~w783;
assign w787 = ~w784 & ~w785;
assign w788 = w786 & w787;
assign w789 = w781 & ~w788;
assign w790 = (~w779 & w777) | (~w779 & w9657) | (w777 & w9657);
assign w791 = ~w789 & w790;
assign w792 = pi1544 & w769;
assign w793 = pi1592 & w773;
assign w794 = pi1568 & w767;
assign w795 = pi1718 & w771;
assign w796 = ~w792 & ~w793;
assign w797 = ~w794 & ~w795;
assign w798 = w796 & w797;
assign w799 = ~pi0243 & w778;
assign w800 = pi1127 & w769;
assign w801 = pi1726 & w771;
assign w802 = pi1112 & w767;
assign w803 = pi1066 & w773;
assign w804 = ~w800 & ~w801;
assign w805 = ~w802 & ~w803;
assign w806 = w804 & w805;
assign w807 = w781 & ~w806;
assign w808 = (~w799 & w798) | (~w799 & w9658) | (w798 & w9658);
assign w809 = ~w807 & w808;
assign w810 = w629 & w9659;
assign w811 = pi1130 & ~pi1183;
assign w812 = w810 & w811;
assign w813 = pi0217 & pi0225;
assign w814 = pi1287 & w813;
assign w815 = ~pi0217 & pi0225;
assign w816 = pi1623 & w815;
assign w817 = pi0217 & ~pi0225;
assign w818 = pi1253 & w817;
assign w819 = ~pi0217 & ~pi0225;
assign w820 = pi1833 & w819;
assign w821 = ~w814 & ~w816;
assign w822 = ~w818 & ~w820;
assign w823 = w821 & w822;
assign w824 = (pi1164 & ~w629) | (pi1164 & w9660) | (~w629 & w9660);
assign w825 = ~pi0244 & w824;
assign w826 = ~pi1130 & pi1183;
assign w827 = w810 & w826;
assign w828 = pi1303 & w813;
assign w829 = pi1048 & w817;
assign w830 = pi1008 & w819;
assign w831 = pi1114 & w815;
assign w832 = ~w828 & ~w829;
assign w833 = ~w830 & ~w831;
assign w834 = w832 & w833;
assign w835 = w827 & ~w834;
assign w836 = (~w825 & w823) | (~w825 & w9661) | (w823 & w9661);
assign w837 = ~w835 & w836;
assign w838 = pi1753 & w819;
assign w839 = pi1281 & w817;
assign w840 = pi1064 & w813;
assign w841 = pi1109 & w815;
assign w842 = ~w838 & ~w839;
assign w843 = ~w840 & ~w841;
assign w844 = w842 & w843;
assign w845 = ~pi0245 & w824;
assign w846 = pi0999 & w819;
assign w847 = pi1649 & w815;
assign w848 = pi1295 & w813;
assign w849 = pi1271 & w817;
assign w850 = ~w846 & ~w847;
assign w851 = ~w848 & ~w849;
assign w852 = w850 & w851;
assign w853 = w812 & ~w852;
assign w854 = (~w845 & w844) | (~w845 & w9662) | (w844 & w9662);
assign w855 = ~w853 & w854;
assign w856 = w621 & w9663;
assign w857 = pi1832 & ~pi1840;
assign w858 = w856 & w857;
assign w859 = pi0216 & ~pi0224;
assign w860 = pi1664 & w859;
assign w861 = ~pi0216 & pi0224;
assign w862 = pi1627 & w861;
assign w863 = pi0216 & pi0224;
assign w864 = pi1257 & w863;
assign w865 = ~pi0216 & ~pi0224;
assign w866 = pi1804 & w865;
assign w867 = ~w860 & ~w862;
assign w868 = ~w864 & ~w866;
assign w869 = w867 & w868;
assign w870 = (pi1838 & ~w621) | (pi1838 & w9664) | (~w621 & w9664);
assign w871 = ~pi0246 & w870;
assign w872 = ~pi1832 & pi1840;
assign w873 = w856 & w872;
assign w874 = pi0995 & w865;
assign w875 = pi1609 & w861;
assign w876 = pi1638 & w859;
assign w877 = pi1231 & w863;
assign w878 = ~w874 & ~w875;
assign w879 = ~w876 & ~w877;
assign w880 = w878 & w879;
assign w881 = w873 & ~w880;
assign w882 = (~w871 & w869) | (~w871 & w9665) | (w869 & w9665);
assign w883 = ~w881 & w882;
assign w884 = pi1051 & w861;
assign w885 = pi1828 & w859;
assign w886 = pi1798 & w865;
assign w887 = pi1098 & w863;
assign w888 = ~w884 & ~w885;
assign w889 = ~w886 & ~w887;
assign w890 = w888 & w889;
assign w891 = ~pi0247 & w870;
assign w892 = pi1617 & w861;
assign w893 = pi1244 & w863;
assign w894 = pi1831 & w865;
assign w895 = pi1652 & w859;
assign w896 = ~w892 & ~w893;
assign w897 = ~w894 & ~w895;
assign w898 = w896 & w897;
assign w899 = w873 & ~w898;
assign w900 = (~w891 & w890) | (~w891 & w9666) | (w890 & w9666);
assign w901 = ~w899 & w900;
assign w902 = ~pi0248 & ~pi0861;
assign w903 = ~w686 & ~w902;
assign w904 = ~pi0249 & ~pi0862;
assign w905 = ~w686 & ~w904;
assign w906 = ~pi0250 & ~pi0863;
assign w907 = ~w686 & ~w906;
assign w908 = ~pi0251 & ~pi0864;
assign w909 = ~w686 & ~w908;
assign w910 = ~pi0252 & w732;
assign w911 = ~w731 & w735;
assign w912 = ~w910 & ~w911;
assign w913 = ~pi0253 & w732;
assign w914 = w735 & ~w752;
assign w915 = ~w913 & ~w914;
assign w916 = ~pi0254 & w778;
assign w917 = ~w777 & w781;
assign w918 = ~w916 & ~w917;
assign w919 = ~pi0255 & w778;
assign w920 = w781 & ~w798;
assign w921 = ~w919 & ~w920;
assign w922 = ~pi0256 & w824;
assign w923 = ~w823 & w827;
assign w924 = ~w922 & ~w923;
assign w925 = w858 & ~w880;
assign w926 = ~pi0257 & w870;
assign w927 = ~w925 & ~w926;
assign w928 = ~pi0258 & w824;
assign w929 = w827 & ~w852;
assign w930 = ~w928 & ~w929;
assign w931 = w858 & ~w898;
assign w932 = ~pi0259 & w870;
assign w933 = ~w931 & ~w932;
assign w934 = w624 & w856;
assign w935 = pi0260 & pi1838;
assign w936 = (w935 & ~w622) | (w935 & w9667) | (~w622 & w9667);
assign w937 = ~w934 & ~w936;
assign w938 = w632 & w810;
assign w939 = pi0261 & pi1164;
assign w940 = (w939 & ~w630) | (w939 & w9668) | (~w630 & w9668);
assign w941 = ~w938 & ~w940;
assign w942 = (~pi0262 & ~w638) | (~pi0262 & w9669) | (~w638 & w9669);
assign w943 = w638 & w9670;
assign w944 = pi1176 & ~w942;
assign w945 = ~w943 & w944;
assign w946 = (~pi0263 & ~w646) | (~pi0263 & w9671) | (~w646 & w9671);
assign w947 = w646 & w9672;
assign w948 = pi1839 & ~w946;
assign w949 = ~w947 & w948;
assign w950 = pi1176 & w943;
assign w951 = pi1522 & w725;
assign w952 = pi1498 & w727;
assign w953 = pi0977 & w721;
assign w954 = pi1474 & w723;
assign w955 = ~w951 & ~w952;
assign w956 = ~w953 & ~w954;
assign w957 = w955 & w956;
assign w958 = w950 & ~w957;
assign w959 = ~pi0264 & w732;
assign w960 = pi1512 & w725;
assign w961 = pi1463 & w723;
assign w962 = pi1081 & w721;
assign w963 = pi1488 & w727;
assign w964 = ~w960 & ~w961;
assign w965 = ~w962 & ~w963;
assign w966 = w964 & w965;
assign w967 = w640 & w718;
assign w968 = pi1713 & w721;
assign w969 = pi1774 & w727;
assign w970 = pi1794 & w723;
assign w971 = pi1124 & w725;
assign w972 = ~w968 & ~w969;
assign w973 = ~w970 & ~w971;
assign w974 = w972 & w973;
assign w975 = w967 & ~w974;
assign w976 = pi1511 & w725;
assign w977 = pi1487 & w727;
assign w978 = pi1462 & w723;
assign w979 = pi1699 & w721;
assign w980 = ~w976 & ~w977;
assign w981 = ~w978 & ~w979;
assign w982 = w980 & w981;
assign w983 = w720 & ~w982;
assign w984 = (~w959 & w966) | (~w959 & w9673) | (w966 & w9673);
assign w985 = ~w975 & ~w983;
assign w986 = w984 & w985;
assign w987 = ~w958 & w986;
assign w988 = pi1499 & w727;
assign w989 = pi1475 & w723;
assign w990 = pi1523 & w725;
assign w991 = pi1708 & w721;
assign w992 = ~w988 & ~w989;
assign w993 = ~w990 & ~w991;
assign w994 = w992 & w993;
assign w995 = w950 & ~w994;
assign w996 = ~pi0265 & w732;
assign w997 = pi1533 & w725;
assign w998 = pi0981 & w721;
assign w999 = pi1509 & w727;
assign w1000 = pi1485 & w723;
assign w1001 = ~w997 & ~w998;
assign w1002 = ~w999 & ~w1000;
assign w1003 = w1001 & w1002;
assign w1004 = pi1464 & w723;
assign w1005 = pi1513 & w725;
assign w1006 = pi1489 & w727;
assign w1007 = pi0972 & w721;
assign w1008 = ~w1004 & ~w1005;
assign w1009 = ~w1006 & ~w1007;
assign w1010 = w1008 & w1009;
assign w1011 = w735 & ~w1010;
assign w1012 = pi1787 & w727;
assign w1013 = pi1802 & w723;
assign w1014 = pi1700 & w721;
assign w1015 = pi1773 & w725;
assign w1016 = ~w1012 & ~w1013;
assign w1017 = ~w1014 & ~w1015;
assign w1018 = w1016 & w1017;
assign w1019 = w720 & ~w1018;
assign w1020 = (~w996 & w1003) | (~w996 & w9674) | (w1003 & w9674);
assign w1021 = ~w1011 & ~w1019;
assign w1022 = w1020 & w1021;
assign w1023 = ~w995 & w1022;
assign w1024 = pi1791 & w723;
assign w1025 = pi1780 & w727;
assign w1026 = pi1706 & w721;
assign w1027 = pi1763 & w725;
assign w1028 = ~w1024 & ~w1025;
assign w1029 = ~w1026 & ~w1027;
assign w1030 = w1028 & w1029;
assign w1031 = w950 & ~w1030;
assign w1032 = ~pi0266 & w732;
assign w1033 = pi1465 & w723;
assign w1034 = pi1514 & w725;
assign w1035 = pi1490 & w727;
assign w1036 = pi0973 & w721;
assign w1037 = ~w1033 & ~w1034;
assign w1038 = ~w1035 & ~w1036;
assign w1039 = w1037 & w1038;
assign w1040 = w735 & ~w1039;
assign w1041 = w720 & ~w966;
assign w1042 = (~w1032 & w982) | (~w1032 & w9675) | (w982 & w9675);
assign w1043 = ~w1040 & ~w1041;
assign w1044 = w1042 & w1043;
assign w1045 = ~w1031 & w1044;
assign w1046 = pi1524 & w725;
assign w1047 = pi1707 & w721;
assign w1048 = pi1476 & w723;
assign w1049 = pi1500 & w727;
assign w1050 = ~w1046 & ~w1047;
assign w1051 = ~w1048 & ~w1049;
assign w1052 = w1050 & w1051;
assign w1053 = w950 & ~w1052;
assign w1054 = ~pi0267 & w732;
assign w1055 = pi1785 & w723;
assign w1056 = pi1784 & w727;
assign w1057 = pi1701 & w721;
assign w1058 = pi1765 & w725;
assign w1059 = ~w1055 & ~w1056;
assign w1060 = ~w1057 & ~w1058;
assign w1061 = w1059 & w1060;
assign w1062 = w735 & ~w1061;
assign w1063 = w720 & ~w1010;
assign w1064 = (~w1054 & w1018) | (~w1054 & w9676) | (w1018 & w9676);
assign w1065 = ~w1062 & ~w1063;
assign w1066 = w1064 & w1065;
assign w1067 = ~w1053 & w1066;
assign w1068 = pi0976 & w721;
assign w1069 = pi1764 & w725;
assign w1070 = pi1757 & w727;
assign w1071 = pi1797 & w723;
assign w1072 = ~w1068 & ~w1069;
assign w1073 = ~w1070 & ~w1071;
assign w1074 = w1072 & w1073;
assign w1075 = w950 & ~w1074;
assign w1076 = ~pi0268 & w732;
assign w1077 = pi1507 & w727;
assign w1078 = pi1118 & w721;
assign w1079 = pi1483 & w723;
assign w1080 = pi1531 & w725;
assign w1081 = ~w1077 & ~w1078;
assign w1082 = ~w1079 & ~w1080;
assign w1083 = w1081 & w1082;
assign w1084 = w967 & ~w1083;
assign w1085 = w735 & ~w982;
assign w1086 = (~w1076 & w974) | (~w1076 & w9677) | (w974 & w9677);
assign w1087 = ~w1084 & ~w1085;
assign w1088 = w1086 & w1087;
assign w1089 = ~w1075 & w1088;
assign w1090 = pi1473 & w723;
assign w1091 = pi1136 & w721;
assign w1092 = pi1497 & w727;
assign w1093 = pi1521 & w725;
assign w1094 = ~w1090 & ~w1091;
assign w1095 = ~w1092 & ~w1093;
assign w1096 = w1094 & w1095;
assign w1097 = w950 & ~w1096;
assign w1098 = ~pi0269 & w732;
assign w1099 = pi1484 & w723;
assign w1100 = pi1508 & w727;
assign w1101 = pi1532 & w725;
assign w1102 = pi0980 & w721;
assign w1103 = ~w1099 & ~w1100;
assign w1104 = ~w1101 & ~w1102;
assign w1105 = w1103 & w1104;
assign w1106 = w720 & ~w1003;
assign w1107 = w735 & ~w1018;
assign w1108 = (~w1098 & w1105) | (~w1098 & w9678) | (w1105 & w9678);
assign w1109 = ~w1106 & ~w1107;
assign w1110 = w1108 & w1109;
assign w1111 = ~w1097 & w1110;
assign w1112 = pi1117 & w721;
assign w1113 = pi1479 & w723;
assign w1114 = pi1527 & w725;
assign w1115 = pi1503 & w727;
assign w1116 = ~w1112 & ~w1113;
assign w1117 = ~w1114 & ~w1115;
assign w1118 = w1116 & w1117;
assign w1119 = w950 & ~w1118;
assign w1120 = ~pi0270 & w732;
assign w1121 = pi1703 & w721;
assign w1122 = pi1493 & w727;
assign w1123 = pi1517 & w725;
assign w1124 = pi1468 & w723;
assign w1125 = ~w1121 & ~w1122;
assign w1126 = ~w1123 & ~w1124;
assign w1127 = w1125 & w1126;
assign w1128 = pi0974 & w721;
assign w1129 = pi1466 & w723;
assign w1130 = pi1515 & w725;
assign w1131 = pi1491 & w727;
assign w1132 = ~w1128 & ~w1129;
assign w1133 = ~w1130 & ~w1131;
assign w1134 = w1132 & w1133;
assign w1135 = w720 & ~w1134;
assign w1136 = w967 & ~w1039;
assign w1137 = (~w1120 & w1127) | (~w1120 & w9679) | (w1127 & w9679);
assign w1138 = ~w1135 & ~w1136;
assign w1139 = w1137 & w1138;
assign w1140 = ~w1119 & w1139;
assign w1141 = pi1528 & w725;
assign w1142 = pi1504 & w727;
assign w1143 = pi1480 & w723;
assign w1144 = pi0978 & w721;
assign w1145 = ~w1141 & ~w1142;
assign w1146 = ~w1143 & ~w1144;
assign w1147 = w1145 & w1146;
assign w1148 = w950 & ~w1147;
assign w1149 = ~pi0271 & w732;
assign w1150 = pi1786 & w727;
assign w1151 = pi1767 & w725;
assign w1152 = pi0975 & w721;
assign w1153 = pi1469 & w723;
assign w1154 = ~w1150 & ~w1151;
assign w1155 = ~w1152 & ~w1153;
assign w1156 = w1154 & w1155;
assign w1157 = pi1447 & w721;
assign w1158 = pi1467 & w723;
assign w1159 = pi1492 & w727;
assign w1160 = pi1516 & w725;
assign w1161 = ~w1157 & ~w1158;
assign w1162 = ~w1159 & ~w1160;
assign w1163 = w1161 & w1162;
assign w1164 = w720 & ~w1163;
assign w1165 = w967 & ~w1061;
assign w1166 = (~w1149 & w1156) | (~w1149 & w9680) | (w1156 & w9680);
assign w1167 = ~w1164 & ~w1165;
assign w1168 = w1166 & w1167;
assign w1169 = ~w1148 & w1168;
assign w1170 = pi1477 & w723;
assign w1171 = pi1501 & w727;
assign w1172 = pi1122 & w721;
assign w1173 = pi1525 & w725;
assign w1174 = ~w1170 & ~w1171;
assign w1175 = ~w1172 & ~w1173;
assign w1176 = w1174 & w1175;
assign w1177 = w950 & ~w1176;
assign w1178 = ~pi0272 & w732;
assign w1179 = ~w966 & w967;
assign w1180 = w735 & ~w1134;
assign w1181 = (~w1178 & w1039) | (~w1178 & w9681) | (w1039 & w9681);
assign w1182 = ~w1179 & ~w1180;
assign w1183 = w1181 & w1182;
assign w1184 = ~w1177 & w1183;
assign w1185 = pi1502 & w727;
assign w1186 = pi1526 & w725;
assign w1187 = pi1710 & w721;
assign w1188 = pi1478 & w723;
assign w1189 = ~w1185 & ~w1186;
assign w1190 = ~w1187 & ~w1188;
assign w1191 = w1189 & w1190;
assign w1192 = w950 & ~w1191;
assign w1193 = ~pi0273 & w732;
assign w1194 = w967 & ~w1010;
assign w1195 = w720 & ~w1061;
assign w1196 = (~w1193 & w1163) | (~w1193 & w9682) | (w1163 & w9682);
assign w1197 = ~w1194 & ~w1195;
assign w1198 = w1196 & w1197;
assign w1199 = ~w1192 & w1198;
assign w1200 = pi0979 & w721;
assign w1201 = pi1759 & w725;
assign w1202 = pi1772 & w727;
assign w1203 = pi1793 & w723;
assign w1204 = ~w1200 & ~w1201;
assign w1205 = ~w1202 & ~w1203;
assign w1206 = w1204 & w1205;
assign w1207 = ~pi0274 & w732;
assign w1208 = w720 & ~w742;
assign w1209 = ~w731 & w967;
assign w1210 = w950 & ~w1134;
assign w1211 = (~w1207 & w1206) | (~w1207 & w9683) | (w1206 & w9683);
assign w1212 = ~w1208 & ~w1209;
assign w1213 = w1211 & w1212;
assign w1214 = ~w1210 & w1213;
assign w1215 = ~pi0275 & w732;
assign w1216 = pi1530 & w725;
assign w1217 = pi1712 & w721;
assign w1218 = pi1506 & w727;
assign w1219 = pi1482 & w723;
assign w1220 = ~w1216 & ~w1217;
assign w1221 = ~w1218 & ~w1219;
assign w1222 = w1220 & w1221;
assign w1223 = w735 & ~w1222;
assign w1224 = ~w752 & w967;
assign w1225 = w950 & ~w1163;
assign w1226 = (~w1215 & w760) | (~w1215 & w9684) | (w760 & w9684);
assign w1227 = ~w1223 & ~w1224;
assign w1228 = w1226 & w1227;
assign w1229 = ~w1225 & w1228;
assign w1230 = w720 & ~w1206;
assign w1231 = w950 & ~w1127;
assign w1232 = ~pi0276 & w732;
assign w1233 = w735 & ~w1083;
assign w1234 = (~w1232 & w742) | (~w1232 & w9685) | (w742 & w9685);
assign w1235 = ~w1230 & ~w1233;
assign w1236 = w1234 & w1235;
assign w1237 = ~w1231 & w1236;
assign w1238 = w720 & ~w1222;
assign w1239 = w950 & ~w1156;
assign w1240 = ~pi0277 & w732;
assign w1241 = w735 & ~w1105;
assign w1242 = (~w1240 & w760) | (~w1240 & w9686) | (w760 & w9686);
assign w1243 = ~w1238 & ~w1241;
assign w1244 = w1242 & w1243;
assign w1245 = ~w1239 & w1244;
assign w1246 = pi1519 & w725;
assign w1247 = pi1471 & w723;
assign w1248 = pi1495 & w727;
assign w1249 = pi1594 & w721;
assign w1250 = ~w1246 & ~w1247;
assign w1251 = ~w1248 & ~w1249;
assign w1252 = w1250 & w1251;
assign w1253 = w950 & ~w1252;
assign w1254 = ~pi0278 & w732;
assign w1255 = w735 & ~w974;
assign w1256 = w967 & ~w1206;
assign w1257 = (~w1254 & w1083) | (~w1254 & w9687) | (w1083 & w9687);
assign w1258 = ~w1255 & ~w1256;
assign w1259 = w1257 & w1258;
assign w1260 = ~w1253 & w1259;
assign w1261 = pi1472 & w723;
assign w1262 = pi1520 & w725;
assign w1263 = pi1705 & w721;
assign w1264 = pi1496 & w727;
assign w1265 = ~w1261 & ~w1262;
assign w1266 = ~w1263 & ~w1264;
assign w1267 = w1265 & w1266;
assign w1268 = w950 & ~w1267;
assign w1269 = ~pi0279 & w732;
assign w1270 = w720 & ~w1105;
assign w1271 = w735 & ~w1003;
assign w1272 = (~w1269 & w1222) | (~w1269 & w9688) | (w1222 & w9688);
assign w1273 = ~w1270 & ~w1271;
assign w1274 = w1272 & w1273;
assign w1275 = ~w1268 & w1274;
assign w1276 = pi1839 & w947;
assign w1277 = pi0986 & w771;
assign w1278 = pi1595 & w773;
assign w1279 = pi1570 & w767;
assign w1280 = pi1546 & w769;
assign w1281 = ~w1277 & ~w1278;
assign w1282 = ~w1279 & ~w1280;
assign w1283 = w1281 & w1282;
assign w1284 = w1276 & ~w1283;
assign w1285 = ~pi0280 & w778;
assign w1286 = w648 & w764;
assign w1287 = pi1581 & w767;
assign w1288 = pi1557 & w769;
assign w1289 = pi1062 & w771;
assign w1290 = pi1606 & w773;
assign w1291 = ~w1287 & ~w1288;
assign w1292 = ~w1289 & ~w1290;
assign w1293 = w1291 & w1292;
assign w1294 = pi1728 & w771;
assign w1295 = pi1558 & w769;
assign w1296 = pi1607 & w773;
assign w1297 = pi1582 & w767;
assign w1298 = ~w1294 & ~w1295;
assign w1299 = ~w1296 & ~w1297;
assign w1300 = w1298 & w1299;
assign w1301 = w766 & ~w1300;
assign w1302 = pi1714 & w771;
assign w1303 = pi1120 & w767;
assign w1304 = pi1107 & w773;
assign w1305 = pi1755 & w769;
assign w1306 = ~w1302 & ~w1303;
assign w1307 = ~w1304 & ~w1305;
assign w1308 = w1306 & w1307;
assign w1309 = w781 & ~w1308;
assign w1310 = (~w1285 & w1293) | (~w1285 & w9689) | (w1293 & w9689);
assign w1311 = ~w1301 & ~w1309;
assign w1312 = w1310 & w1311;
assign w1313 = ~w1284 & w1312;
assign w1314 = pi1073 & w771;
assign w1315 = pi1596 & w773;
assign w1316 = pi1547 & w769;
assign w1317 = pi1571 & w767;
assign w1318 = ~w1314 & ~w1315;
assign w1319 = ~w1316 & ~w1317;
assign w1320 = w1318 & w1319;
assign w1321 = w1276 & ~w1320;
assign w1322 = ~pi0281 & w778;
assign w1323 = pi1608 & w773;
assign w1324 = pi0991 & w771;
assign w1325 = pi1583 & w767;
assign w1326 = pi1559 & w769;
assign w1327 = ~w1323 & ~w1324;
assign w1328 = ~w1325 & ~w1326;
assign w1329 = w1327 & w1328;
assign w1330 = pi1083 & w773;
assign w1331 = pi0990 & w771;
assign w1332 = pi1106 & w767;
assign w1333 = pi1123 & w769;
assign w1334 = ~w1330 & ~w1331;
assign w1335 = ~w1332 & ~w1333;
assign w1336 = w1334 & w1335;
assign w1337 = w1286 & ~w1336;
assign w1338 = pi1585 & w773;
assign w1339 = pi1536 & w769;
assign w1340 = pi1715 & w771;
assign w1341 = pi1561 & w767;
assign w1342 = ~w1338 & ~w1339;
assign w1343 = ~w1340 & ~w1341;
assign w1344 = w1342 & w1343;
assign w1345 = w781 & ~w1344;
assign w1346 = (~w1322 & w1329) | (~w1322 & w9690) | (w1329 & w9690);
assign w1347 = ~w1337 & ~w1345;
assign w1348 = w1346 & w1347;
assign w1349 = ~w1321 & w1348;
assign w1350 = pi1572 & w767;
assign w1351 = pi1548 & w769;
assign w1352 = pi0987 & w771;
assign w1353 = pi1597 & w773;
assign w1354 = ~w1350 & ~w1351;
assign w1355 = ~w1352 & ~w1353;
assign w1356 = w1354 & w1355;
assign w1357 = w1276 & ~w1356;
assign w1358 = ~pi0282 & w778;
assign w1359 = pi1562 & w767;
assign w1360 = pi1586 & w773;
assign w1361 = pi1087 & w771;
assign w1362 = pi1537 & w769;
assign w1363 = ~w1359 & ~w1360;
assign w1364 = ~w1361 & ~w1362;
assign w1365 = w1363 & w1364;
assign w1366 = w1286 & ~w1300;
assign w1367 = w766 & ~w1308;
assign w1368 = (~w1358 & w1365) | (~w1358 & w9691) | (w1365 & w9691);
assign w1369 = ~w1366 & ~w1367;
assign w1370 = w1368 & w1369;
assign w1371 = ~w1357 & w1370;
assign w1372 = pi1720 & w771;
assign w1373 = pi1105 & w767;
assign w1374 = pi1063 & w769;
assign w1375 = pi1089 & w773;
assign w1376 = ~w1372 & ~w1373;
assign w1377 = ~w1374 & ~w1375;
assign w1378 = w1376 & w1377;
assign w1379 = w1276 & ~w1378;
assign w1380 = ~pi0283 & w778;
assign w1381 = pi1587 & w773;
assign w1382 = pi1563 & w767;
assign w1383 = pi0982 & w771;
assign w1384 = pi1538 & w769;
assign w1385 = ~w1381 & ~w1382;
assign w1386 = ~w1383 & ~w1384;
assign w1387 = w1385 & w1386;
assign w1388 = w781 & ~w1387;
assign w1389 = w766 & ~w1344;
assign w1390 = (~w1380 & w1329) | (~w1380 & w9692) | (w1329 & w9692);
assign w1391 = ~w1388 & ~w1389;
assign w1392 = w1390 & w1391;
assign w1393 = ~w1379 & w1392;
assign w1394 = pi1549 & w769;
assign w1395 = pi1598 & w773;
assign w1396 = pi1723 & w771;
assign w1397 = pi1573 & w767;
assign w1398 = ~w1394 & ~w1395;
assign w1399 = ~w1396 & ~w1397;
assign w1400 = w1398 & w1399;
assign w1401 = w1276 & ~w1400;
assign w1402 = ~pi0284 & w778;
assign w1403 = pi1391 & w769;
assign w1404 = pi1119 & w767;
assign w1405 = pi1088 & w773;
assign w1406 = pi0983 & w771;
assign w1407 = ~w1403 & ~w1404;
assign w1408 = ~w1405 & ~w1406;
assign w1409 = w1407 & w1408;
assign w1410 = w781 & ~w1409;
assign w1411 = w1286 & ~w1308;
assign w1412 = (~w1402 & w1365) | (~w1402 & w9693) | (w1365 & w9693);
assign w1413 = ~w1410 & ~w1411;
assign w1414 = w1412 & w1413;
assign w1415 = ~w1401 & w1414;
assign w1416 = pi1135 & w769;
assign w1417 = pi1090 & w773;
assign w1418 = pi1725 & w771;
assign w1419 = pi1113 & w767;
assign w1420 = ~w1416 & ~w1417;
assign w1421 = ~w1418 & ~w1419;
assign w1422 = w1420 & w1421;
assign w1423 = w1276 & ~w1422;
assign w1424 = ~pi0285 & w778;
assign w1425 = pi1716 & w771;
assign w1426 = pi1588 & w773;
assign w1427 = pi1539 & w769;
assign w1428 = pi1564 & w767;
assign w1429 = ~w1425 & ~w1426;
assign w1430 = ~w1427 & ~w1428;
assign w1431 = w1429 & w1430;
assign w1432 = w1286 & ~w1387;
assign w1433 = pi1101 & w771;
assign w1434 = pi1541 & w769;
assign w1435 = pi1590 & w773;
assign w1436 = pi1566 & w767;
assign w1437 = ~w1433 & ~w1434;
assign w1438 = ~w1435 & ~w1436;
assign w1439 = w1437 & w1438;
assign w1440 = w781 & ~w1439;
assign w1441 = (~w1424 & w1431) | (~w1424 & w9694) | (w1431 & w9694);
assign w1442 = ~w1432 & ~w1440;
assign w1443 = w1441 & w1442;
assign w1444 = ~w1423 & w1443;
assign w1445 = pi1721 & w771;
assign w1446 = pi1550 & w769;
assign w1447 = pi1599 & w773;
assign w1448 = pi1574 & w767;
assign w1449 = ~w1445 & ~w1446;
assign w1450 = ~w1447 & ~w1448;
assign w1451 = w1449 & w1450;
assign w1452 = w1276 & ~w1451;
assign w1453 = ~pi0286 & w778;
assign w1454 = w781 & ~w1431;
assign w1455 = w766 & ~w1387;
assign w1456 = (~w1453 & w1344) | (~w1453 & w9695) | (w1344 & w9695);
assign w1457 = ~w1454 & ~w1455;
assign w1458 = w1456 & w1457;
assign w1459 = ~w1452 & w1458;
assign w1460 = pi1578 & w767;
assign w1461 = pi1603 & w773;
assign w1462 = pi1554 & w769;
assign w1463 = pi0988 & w771;
assign w1464 = ~w1460 & ~w1461;
assign w1465 = ~w1462 & ~w1463;
assign w1466 = w1464 & w1465;
assign w1467 = w1276 & ~w1466;
assign w1468 = ~pi0287 & w778;
assign w1469 = pi1591 & w773;
assign w1470 = pi0985 & w771;
assign w1471 = pi1567 & w767;
assign w1472 = pi1543 & w769;
assign w1473 = ~w1469 & ~w1470;
assign w1474 = ~w1471 & ~w1472;
assign w1475 = w1473 & w1474;
assign w1476 = w766 & ~w1439;
assign w1477 = w1286 & ~w1431;
assign w1478 = (~w1468 & w1475) | (~w1468 & w9696) | (w1475 & w9696);
assign w1479 = ~w1476 & ~w1477;
assign w1480 = w1478 & w1479;
assign w1481 = ~w1467 & w1480;
assign w1482 = pi1575 & w767;
assign w1483 = pi1600 & w773;
assign w1484 = pi1722 & w771;
assign w1485 = pi1551 & w769;
assign w1486 = ~w1482 & ~w1483;
assign w1487 = ~w1484 & ~w1485;
assign w1488 = w1486 & w1487;
assign w1489 = w1276 & ~w1488;
assign w1490 = ~pi0288 & w778;
assign w1491 = w1286 & ~w1365;
assign w1492 = pi1565 & w767;
assign w1493 = pi0984 & w771;
assign w1494 = pi1540 & w769;
assign w1495 = pi1589 & w773;
assign w1496 = ~w1492 & ~w1493;
assign w1497 = ~w1494 & ~w1495;
assign w1498 = w1496 & w1497;
assign w1499 = w781 & ~w1498;
assign w1500 = (~w1490 & w1409) | (~w1490 & w9697) | (w1409 & w9697);
assign w1501 = ~w1491 & ~w1499;
assign w1502 = w1500 & w1501;
assign w1503 = ~w1489 & w1502;
assign w1504 = pi1047 & w771;
assign w1505 = pi1602 & w773;
assign w1506 = pi1577 & w767;
assign w1507 = pi1553 & w769;
assign w1508 = ~w1504 & ~w1505;
assign w1509 = ~w1506 & ~w1507;
assign w1510 = w1508 & w1509;
assign w1511 = w1276 & ~w1510;
assign w1512 = ~pi0289 & w778;
assign w1513 = pi1097 & w773;
assign w1514 = pi1116 & w767;
assign w1515 = pi1717 & w771;
assign w1516 = pi1542 & w769;
assign w1517 = ~w1513 & ~w1514;
assign w1518 = ~w1515 & ~w1516;
assign w1519 = w1517 & w1518;
assign w1520 = w766 & ~w1498;
assign w1521 = w1286 & ~w1409;
assign w1522 = (~w1512 & w1519) | (~w1512 & w9698) | (w1519 & w9698);
assign w1523 = ~w1520 & ~w1521;
assign w1524 = w1522 & w1523;
assign w1525 = ~w1511 & w1524;
assign w1526 = ~pi0290 & w778;
assign w1527 = pi1555 & w769;
assign w1528 = pi1604 & w773;
assign w1529 = pi1579 & w767;
assign w1530 = pi0989 & w771;
assign w1531 = ~w1527 & ~w1528;
assign w1532 = ~w1529 & ~w1530;
assign w1533 = w1531 & w1532;
assign w1534 = w781 & ~w1533;
assign w1535 = w766 & ~w788;
assign w1536 = w1276 & ~w1498;
assign w1537 = (~w1526 & w777) | (~w1526 & w9699) | (w777 & w9699);
assign w1538 = ~w1534 & ~w1535;
assign w1539 = w1537 & w1538;
assign w1540 = ~w1536 & w1539;
assign w1541 = ~pi0291 & w778;
assign w1542 = pi1580 & w767;
assign w1543 = pi1556 & w769;
assign w1544 = pi1605 & w773;
assign w1545 = pi1727 & w771;
assign w1546 = ~w1542 & ~w1543;
assign w1547 = ~w1544 & ~w1545;
assign w1548 = w1546 & w1547;
assign w1549 = w781 & ~w1548;
assign w1550 = w766 & ~w806;
assign w1551 = w1276 & ~w1439;
assign w1552 = (~w1541 & w798) | (~w1541 & w9700) | (w798 & w9700);
assign w1553 = ~w1549 & ~w1550;
assign w1554 = w1552 & w1553;
assign w1555 = ~w1551 & w1554;
assign w1556 = w781 & ~w1293;
assign w1557 = w1276 & ~w1519;
assign w1558 = ~pi0292 & w778;
assign w1559 = ~w788 & w1286;
assign w1560 = (~w1558 & w1533) | (~w1558 & w9701) | (w1533 & w9701);
assign w1561 = ~w1556 & ~w1559;
assign w1562 = w1560 & w1561;
assign w1563 = ~w1557 & w1562;
assign w1564 = ~w806 & w1286;
assign w1565 = w1276 & ~w1475;
assign w1566 = ~pi0293 & w778;
assign w1567 = w766 & ~w1548;
assign w1568 = (~w1566 & w1336) | (~w1566 & w9702) | (w1336 & w9702);
assign w1569 = ~w1564 & ~w1567;
assign w1570 = w1568 & w1569;
assign w1571 = ~w1565 & w1570;
assign w1572 = pi1545 & w769;
assign w1573 = pi1015 & w771;
assign w1574 = pi1569 & w767;
assign w1575 = pi1593 & w773;
assign w1576 = ~w1572 & ~w1573;
assign w1577 = ~w1574 & ~w1575;
assign w1578 = w1576 & w1577;
assign w1579 = w1276 & ~w1578;
assign w1580 = ~pi0294 & w778;
assign w1581 = w1286 & ~w1533;
assign w1582 = w781 & ~w1300;
assign w1583 = (~w1580 & w1293) | (~w1580 & w9703) | (w1293 & w9703);
assign w1584 = ~w1581 & ~w1582;
assign w1585 = w1583 & w1584;
assign w1586 = ~w1579 & w1585;
assign w1587 = pi1096 & w773;
assign w1588 = pi1702 & w769;
assign w1589 = pi1115 & w767;
assign w1590 = pi1719 & w771;
assign w1591 = ~w1587 & ~w1588;
assign w1592 = ~w1589 & ~w1590;
assign w1593 = w1591 & w1592;
assign w1594 = w1276 & ~w1593;
assign w1595 = ~pi0295 & w778;
assign w1596 = w1286 & ~w1548;
assign w1597 = w781 & ~w1329;
assign w1598 = (~w1595 & w1336) | (~w1595 & w9704) | (w1336 & w9704);
assign w1599 = ~w1596 & ~w1597;
assign w1600 = w1598 & w1599;
assign w1601 = ~w1594 & w1600;
assign w1602 = pi1729 & w819;
assign w1603 = pi1625 & w815;
assign w1604 = pi1255 & w817;
assign w1605 = pi1288 & w813;
assign w1606 = ~w1602 & ~w1603;
assign w1607 = ~w1604 & ~w1605;
assign w1608 = w1606 & w1607;
assign w1609 = ~pi0296 & w824;
assign w1610 = pi1754 & w819;
assign w1611 = pi1534 & w813;
assign w1612 = pi1248 & w815;
assign w1613 = pi1086 & w817;
assign w1614 = ~w1610 & ~w1611;
assign w1615 = ~w1612 & ~w1613;
assign w1616 = w1614 & w1615;
assign w1617 = w812 & ~w1616;
assign w1618 = pi1243 & w815;
assign w1619 = pi1010 & w819;
assign w1620 = pi1069 & w813;
assign w1621 = pi1284 & w817;
assign w1622 = ~w1618 & ~w1619;
assign w1623 = ~w1620 & ~w1621;
assign w1624 = w1622 & w1623;
assign w1625 = w938 & ~w1624;
assign w1626 = w630 & w9705;
assign w1627 = pi1092 & w817;
assign w1628 = pi1025 & w815;
assign w1629 = pi1740 & w819;
assign w1630 = pi1070 & w813;
assign w1631 = ~w1627 & ~w1628;
assign w1632 = ~w1629 & ~w1630;
assign w1633 = w1631 & w1632;
assign w1634 = w1626 & ~w1633;
assign w1635 = (~w1609 & w1608) | (~w1609 & w9706) | (w1608 & w9706);
assign w1636 = ~w1617 & ~w1625;
assign w1637 = ~w1634 & w1636;
assign w1638 = w1635 & w1637;
assign w1639 = pi1050 & w815;
assign w1640 = pi1099 & w817;
assign w1641 = pi0992 & w819;
assign w1642 = pi1085 & w813;
assign w1643 = ~w1639 & ~w1640;
assign w1644 = ~w1641 & ~w1642;
assign w1645 = w1643 & w1644;
assign w1646 = ~pi0297 & w824;
assign w1647 = pi1286 & w817;
assign w1648 = pi1251 & w815;
assign w1649 = pi1776 & w819;
assign w1650 = pi1308 & w813;
assign w1651 = ~w1647 & ~w1648;
assign w1652 = ~w1649 & ~w1650;
assign w1653 = w1651 & w1652;
assign w1654 = w812 & ~w1653;
assign w1655 = pi1855 & w819;
assign w1656 = pi1307 & w813;
assign w1657 = pi1245 & w815;
assign w1658 = pi1285 & w817;
assign w1659 = ~w1655 & ~w1656;
assign w1660 = ~w1657 & ~w1658;
assign w1661 = w1659 & w1660;
assign w1662 = w938 & ~w1661;
assign w1663 = pi1273 & w817;
assign w1664 = pi1658 & w815;
assign w1665 = pi1807 & w819;
assign w1666 = pi1298 & w813;
assign w1667 = ~w1663 & ~w1664;
assign w1668 = ~w1665 & ~w1666;
assign w1669 = w1667 & w1668;
assign w1670 = w1626 & ~w1669;
assign w1671 = (~w1646 & w1645) | (~w1646 & w9707) | (w1645 & w9707);
assign w1672 = ~w1654 & ~w1662;
assign w1673 = ~w1670 & w1672;
assign w1674 = w1671 & w1673;
assign w1675 = ~pi0298 & w824;
assign w1676 = pi1632 & w815;
assign w1677 = pi1262 & w817;
assign w1678 = pi1058 & w819;
assign w1679 = pi1290 & w813;
assign w1680 = ~w1676 & ~w1677;
assign w1681 = ~w1678 & ~w1679;
assign w1682 = w1680 & w1681;
assign w1683 = w827 & ~w1682;
assign w1684 = w938 & ~w1653;
assign w1685 = pi1309 & w813;
assign w1686 = pi1662 & w815;
assign w1687 = pi1275 & w817;
assign w1688 = pi1745 & w819;
assign w1689 = ~w1685 & ~w1686;
assign w1690 = ~w1687 & ~w1688;
assign w1691 = w1689 & w1690;
assign w1692 = w1626 & ~w1691;
assign w1693 = (~w1675 & w1645) | (~w1675 & w9708) | (w1645 & w9708);
assign w1694 = ~w1683 & ~w1684;
assign w1695 = ~w1692 & w1694;
assign w1696 = w1693 & w1695;
assign w1697 = pi1264 & w817;
assign w1698 = pi1854 & w819;
assign w1699 = pi1291 & w813;
assign w1700 = pi1634 & w815;
assign w1701 = ~w1697 & ~w1698;
assign w1702 = ~w1699 & ~w1700;
assign w1703 = w1701 & w1702;
assign w1704 = ~pi0299 & w824;
assign w1705 = pi1630 & w815;
assign w1706 = pi1289 & w813;
assign w1707 = pi0993 & w819;
assign w1708 = pi1260 & w817;
assign w1709 = ~w1705 & ~w1706;
assign w1710 = ~w1707 & ~w1708;
assign w1711 = w1709 & w1710;
assign w1712 = w812 & ~w1711;
assign w1713 = w938 & ~w1608;
assign w1714 = pi1824 & w815;
assign w1715 = pi1091 & w817;
assign w1716 = pi1300 & w813;
assign w1717 = pi1746 & w819;
assign w1718 = ~w1714 & ~w1715;
assign w1719 = ~w1716 & ~w1717;
assign w1720 = w1718 & w1719;
assign w1721 = w1626 & ~w1720;
assign w1722 = (~w1704 & w1703) | (~w1704 & w9709) | (w1703 & w9709);
assign w1723 = ~w1712 & ~w1713;
assign w1724 = ~w1721 & w1723;
assign w1725 = w1722 & w1724;
assign w1726 = ~pi0300 & w824;
assign w1727 = pi1043 & w815;
assign w1728 = pi0994 & w819;
assign w1729 = pi1266 & w817;
assign w1730 = pi1084 & w813;
assign w1731 = ~w1727 & ~w1728;
assign w1732 = ~w1729 & ~w1730;
assign w1733 = w1731 & w1732;
assign w1734 = w827 & ~w1733;
assign w1735 = w938 & ~w1645;
assign w1736 = pi1276 & w817;
assign w1737 = pi1072 & w813;
assign w1738 = pi1667 & w815;
assign w1739 = pi1005 & w819;
assign w1740 = ~w1736 & ~w1737;
assign w1741 = ~w1738 & ~w1739;
assign w1742 = w1740 & w1741;
assign w1743 = w1626 & ~w1742;
assign w1744 = (~w1726 & w1682) | (~w1726 & w9710) | (w1682 & w9710);
assign w1745 = ~w1734 & ~w1735;
assign w1746 = ~w1743 & w1745;
assign w1747 = w1744 & w1746;
assign w1748 = ~pi0301 & w824;
assign w1749 = pi1292 & w813;
assign w1750 = pi1639 & w815;
assign w1751 = pi1268 & w817;
assign w1752 = pi1031 & w819;
assign w1753 = ~w1749 & ~w1750;
assign w1754 = ~w1751 & ~w1752;
assign w1755 = w1753 & w1754;
assign w1756 = w827 & ~w1755;
assign w1757 = w938 & ~w1711;
assign w1758 = pi1225 & w815;
assign w1759 = pi1747 & w819;
assign w1760 = pi1277 & w817;
assign w1761 = pi1301 & w813;
assign w1762 = ~w1758 & ~w1759;
assign w1763 = ~w1760 & ~w1761;
assign w1764 = w1762 & w1763;
assign w1765 = w1626 & ~w1764;
assign w1766 = (~w1748 & w1703) | (~w1748 & w9711) | (w1703 & w9711);
assign w1767 = ~w1756 & ~w1757;
assign w1768 = ~w1765 & w1767;
assign w1769 = w1766 & w1768;
assign w1770 = ~pi0302 & w824;
assign w1771 = pi1269 & w817;
assign w1772 = pi1293 & w813;
assign w1773 = pi1642 & w815;
assign w1774 = pi1013 & w819;
assign w1775 = ~w1771 & ~w1772;
assign w1776 = ~w1773 & ~w1774;
assign w1777 = w1775 & w1776;
assign w1778 = w827 & ~w1777;
assign w1779 = w938 & ~w1682;
assign w1780 = pi1278 & w817;
assign w1781 = pi1227 & w815;
assign w1782 = pi1302 & w813;
assign w1783 = pi1009 & w819;
assign w1784 = ~w1780 & ~w1781;
assign w1785 = ~w1782 & ~w1783;
assign w1786 = w1784 & w1785;
assign w1787 = w1626 & ~w1786;
assign w1788 = (~w1770 & w1733) | (~w1770 & w9712) | (w1733 & w9712);
assign w1789 = ~w1778 & ~w1779;
assign w1790 = ~w1787 & w1789;
assign w1791 = w1788 & w1790;
assign w1792 = pi1093 & w817;
assign w1793 = pi1294 & w813;
assign w1794 = pi1732 & w819;
assign w1795 = pi1644 & w815;
assign w1796 = ~w1792 & ~w1793;
assign w1797 = ~w1794 & ~w1795;
assign w1798 = w1796 & w1797;
assign w1799 = ~pi0303 & w824;
assign w1800 = w812 & ~w1755;
assign w1801 = pi1232 & w815;
assign w1802 = pi1279 & w817;
assign w1803 = pi1752 & w819;
assign w1804 = pi1071 & w813;
assign w1805 = ~w1801 & ~w1802;
assign w1806 = ~w1803 & ~w1804;
assign w1807 = w1805 & w1806;
assign w1808 = w1626 & ~w1807;
assign w1809 = w938 & ~w1703;
assign w1810 = (~w1799 & w1798) | (~w1799 & w9713) | (w1798 & w9713);
assign w1811 = ~w1800 & ~w1808;
assign w1812 = ~w1809 & w1811;
assign w1813 = w1810 & w1812;
assign w1814 = pi1121 & w859;
assign w1815 = pi1034 & w861;
assign w1816 = pi1095 & w863;
assign w1817 = pi1750 & w865;
assign w1818 = ~w1814 & ~w1815;
assign w1819 = ~w1816 & ~w1817;
assign w1820 = w1818 & w1819;
assign w1821 = ~pi0304 & w870;
assign w1822 = pi1082 & w861;
assign w1823 = pi1730 & w865;
assign w1824 = pi1111 & w863;
assign w1825 = pi1640 & w859;
assign w1826 = ~w1822 & ~w1823;
assign w1827 = ~w1824 & ~w1825;
assign w1828 = w1826 & w1827;
assign w1829 = w858 & ~w1828;
assign w1830 = pi1749 & w865;
assign w1831 = pi1229 & w859;
assign w1832 = pi1636 & w861;
assign w1833 = pi1094 & w863;
assign w1834 = ~w1830 & ~w1831;
assign w1835 = ~w1832 & ~w1833;
assign w1836 = w1834 & w1835;
assign w1837 = w873 & ~w1836;
assign w1838 = w622 & w9714;
assign w1839 = pi1103 & w863;
assign w1840 = pi1619 & w861;
assign w1841 = pi1820 & w865;
assign w1842 = pi1655 & w859;
assign w1843 = ~w1839 & ~w1840;
assign w1844 = ~w1841 & ~w1842;
assign w1845 = w1843 & w1844;
assign w1846 = w1838 & ~w1845;
assign w1847 = (~w1821 & w1820) | (~w1821 & w9715) | (w1820 & w9715);
assign w1848 = ~w1829 & ~w1837;
assign w1849 = ~w1846 & w1848;
assign w1850 = w1847 & w1849;
assign w1851 = pi1734 & w819;
assign w1852 = pi1038 & w815;
assign w1853 = pi1074 & w813;
assign w1854 = pi1270 & w817;
assign w1855 = ~w1851 & ~w1852;
assign w1856 = ~w1853 & ~w1854;
assign w1857 = w1855 & w1856;
assign w1858 = ~pi0305 & w824;
assign w1859 = w938 & ~w1733;
assign w1860 = pi1304 & w813;
assign w1861 = pi1872 & w819;
assign w1862 = pi1280 & w817;
assign w1863 = pi1234 & w815;
assign w1864 = ~w1860 & ~w1861;
assign w1865 = ~w1862 & ~w1863;
assign w1866 = w1864 & w1865;
assign w1867 = w1626 & ~w1866;
assign w1868 = w812 & ~w1777;
assign w1869 = (~w1858 & w1857) | (~w1858 & w9716) | (w1857 & w9716);
assign w1870 = ~w1859 & ~w1867;
assign w1871 = ~w1868 & w1870;
assign w1872 = w1869 & w1871;
assign w1873 = pi1751 & w865;
assign w1874 = pi1637 & w861;
assign w1875 = pi1230 & w859;
assign w1876 = pi1267 & w863;
assign w1877 = ~w1873 & ~w1874;
assign w1878 = ~w1875 & ~w1876;
assign w1879 = w1877 & w1878;
assign w1880 = ~pi0306 & w870;
assign w1881 = pi0996 & w865;
assign w1882 = pi1641 & w859;
assign w1883 = pi1610 & w861;
assign w1884 = pi1233 & w863;
assign w1885 = ~w1881 & ~w1882;
assign w1886 = ~w1883 & ~w1884;
assign w1887 = w1885 & w1886;
assign w1888 = w858 & ~w1887;
assign w1889 = pi1748 & w865;
assign w1890 = pi1635 & w861;
assign w1891 = pi1265 & w863;
assign w1892 = pi1228 & w859;
assign w1893 = ~w1889 & ~w1890;
assign w1894 = ~w1891 & ~w1892;
assign w1895 = w1893 & w1894;
assign w1896 = w934 & ~w1895;
assign w1897 = pi1656 & w859;
assign w1898 = pi1249 & w863;
assign w1899 = pi1620 & w861;
assign w1900 = pi1741 & w865;
assign w1901 = ~w1897 & ~w1898;
assign w1902 = ~w1899 & ~w1900;
assign w1903 = w1901 & w1902;
assign w1904 = w1838 & ~w1903;
assign w1905 = (~w1880 & w1879) | (~w1880 & w9717) | (w1879 & w9717);
assign w1906 = ~w1888 & ~w1896;
assign w1907 = ~w1904 & w1906;
assign w1908 = w1905 & w1907;
assign w1909 = ~pi0307 & w870;
assign w1910 = w873 & ~w1828;
assign w1911 = pi1235 & w863;
assign w1912 = pi1611 & w861;
assign w1913 = pi1643 & w859;
assign w1914 = pi0997 & w865;
assign w1915 = ~w1911 & ~w1912;
assign w1916 = ~w1913 & ~w1914;
assign w1917 = w1915 & w1916;
assign w1918 = w858 & ~w1917;
assign w1919 = pi1742 & w865;
assign w1920 = pi1657 & w859;
assign w1921 = pi1250 & w863;
assign w1922 = pi1621 & w861;
assign w1923 = ~w1919 & ~w1920;
assign w1924 = ~w1921 & ~w1922;
assign w1925 = w1923 & w1924;
assign w1926 = w1838 & ~w1925;
assign w1927 = (~w1909 & w1836) | (~w1909 & w9718) | (w1836 & w9718);
assign w1928 = ~w1910 & ~w1918;
assign w1929 = ~w1926 & w1928;
assign w1930 = w1927 & w1929;
assign w1931 = ~pi0308 & w824;
assign w1932 = w812 & ~w1608;
assign w1933 = w938 & ~w1616;
assign w1934 = pi1660 & w815;
assign w1935 = pi1274 & w817;
assign w1936 = pi1299 & w813;
assign w1937 = pi1744 & w819;
assign w1938 = ~w1934 & ~w1935;
assign w1939 = ~w1936 & ~w1937;
assign w1940 = w1938 & w1939;
assign w1941 = w1626 & ~w1940;
assign w1942 = (~w1931 & w1711) | (~w1931 & w9719) | (w1711 & w9719);
assign w1943 = ~w1932 & ~w1933;
assign w1944 = ~w1941 & w1943;
assign w1945 = w1942 & w1944;
assign w1946 = ~pi0309 & w870;
assign w1947 = pi1731 & w865;
assign w1948 = pi1612 & w861;
assign w1949 = pi1037 & w859;
assign w1950 = pi1236 & w863;
assign w1951 = ~w1947 & ~w1948;
assign w1952 = ~w1949 & ~w1950;
assign w1953 = w1951 & w1952;
assign w1954 = w858 & ~w1953;
assign w1955 = w934 & ~w1879;
assign w1956 = pi1104 & w863;
assign w1957 = pi1016 & w859;
assign w1958 = pi1059 & w861;
assign w1959 = pi1743 & w865;
assign w1960 = ~w1956 & ~w1957;
assign w1961 = ~w1958 & ~w1959;
assign w1962 = w1960 & w1961;
assign w1963 = w1838 & ~w1962;
assign w1964 = (~w1946 & w1887) | (~w1946 & w9720) | (w1887 & w9720);
assign w1965 = ~w1954 & ~w1955;
assign w1966 = ~w1963 & w1965;
assign w1967 = w1964 & w1966;
assign w1968 = pi1645 & w859;
assign w1969 = pi1238 & w863;
assign w1970 = pi1733 & w865;
assign w1971 = pi1067 & w861;
assign w1972 = ~w1968 & ~w1969;
assign w1973 = ~w1970 & ~w1971;
assign w1974 = w1972 & w1973;
assign w1975 = ~pi0310 & w870;
assign w1976 = w934 & ~w1828;
assign w1977 = w873 & ~w1917;
assign w1978 = pi1001 & w865;
assign w1979 = pi1622 & w861;
assign w1980 = pi1252 & w863;
assign w1981 = pi1659 & w859;
assign w1982 = ~w1978 & ~w1979;
assign w1983 = ~w1980 & ~w1981;
assign w1984 = w1982 & w1983;
assign w1985 = w1838 & ~w1984;
assign w1986 = (~w1975 & w1974) | (~w1975 & w9721) | (w1974 & w9721);
assign w1987 = ~w1976 & ~w1977;
assign w1988 = ~w1985 & w1987;
assign w1989 = w1986 & w1988;
assign w1990 = ~pi0311 & w824;
assign w1991 = pi1781 & w819;
assign w1992 = pi1305 & w813;
assign w1993 = pi1237 & w815;
assign w1994 = pi1282 & w817;
assign w1995 = ~w1991 & ~w1992;
assign w1996 = ~w1993 & ~w1994;
assign w1997 = w1995 & w1996;
assign w1998 = w827 & ~w1997;
assign w1999 = ~w823 & w938;
assign w2000 = w812 & ~w834;
assign w2001 = (~w1990 & w1755) | (~w1990 & w9722) | (w1755 & w9722);
assign w2002 = ~w1998 & ~w1999;
assign w2003 = ~w2000 & w2002;
assign w2004 = w2001 & w2003;
assign w2005 = pi1647 & w859;
assign w2006 = pi1800 & w865;
assign w2007 = pi1239 & w863;
assign w2008 = pi1614 & w861;
assign w2009 = ~w2005 & ~w2006;
assign w2010 = ~w2007 & ~w2008;
assign w2011 = w2009 & w2010;
assign w2012 = ~pi0312 & w870;
assign w2013 = w873 & ~w1974;
assign w2014 = w934 & ~w1917;
assign w2015 = pi1057 & w861;
assign w2016 = pi1002 & w865;
assign w2017 = pi1017 & w859;
assign w2018 = pi1100 & w863;
assign w2019 = ~w2015 & ~w2016;
assign w2020 = ~w2017 & ~w2018;
assign w2021 = w2019 & w2020;
assign w2022 = w1838 & ~w2021;
assign w2023 = (~w2012 & w2011) | (~w2012 & w9723) | (w2011 & w9723);
assign w2024 = ~w2013 & ~w2014;
assign w2025 = ~w2022 & w2024;
assign w2026 = w2023 & w2025;
assign w2027 = ~pi0313 & w824;
assign w2028 = ~w834 & w938;
assign w2029 = w827 & ~w1624;
assign w2030 = w1626 & ~w1798;
assign w2031 = (~w2027 & w1997) | (~w2027 & w9724) | (w1997 & w9724);
assign w2032 = ~w2028 & ~w2029;
assign w2033 = ~w2030 & w2032;
assign w2034 = w2031 & w2033;
assign w2035 = pi0998 & w865;
assign w2036 = pi1615 & w861;
assign w2037 = pi1648 & w859;
assign w2038 = pi1240 & w863;
assign w2039 = ~w2035 & ~w2036;
assign w2040 = ~w2037 & ~w2038;
assign w2041 = w2039 & w2040;
assign w2042 = ~pi0314 & w870;
assign w2043 = pi1646 & w859;
assign w2044 = pi1030 & w865;
assign w2045 = pi1110 & w863;
assign w2046 = pi1613 & w861;
assign w2047 = ~w2043 & ~w2044;
assign w2048 = ~w2045 & ~w2046;
assign w2049 = w2047 & w2048;
assign w2050 = w873 & ~w2049;
assign w2051 = w934 & ~w1953;
assign w2052 = pi1256 & w863;
assign w2053 = pi1663 & w859;
assign w2054 = pi1003 & w865;
assign w2055 = pi1626 & w861;
assign w2056 = ~w2052 & ~w2053;
assign w2057 = ~w2054 & ~w2055;
assign w2058 = w2056 & w2057;
assign w2059 = w1838 & ~w2058;
assign w2060 = (~w2042 & w2041) | (~w2042 & w9725) | (w2041 & w9725);
assign w2061 = ~w2050 & ~w2051;
assign w2062 = ~w2059 & w2061;
assign w2063 = w2060 & w2062;
assign w2064 = pi1011 & w819;
assign w2065 = pi1283 & w817;
assign w2066 = pi1306 & w813;
assign w2067 = pi1241 & w815;
assign w2068 = ~w2064 & ~w2065;
assign w2069 = ~w2066 & ~w2067;
assign w2070 = w2068 & w2069;
assign w2071 = ~pi0315 & w824;
assign w2072 = ~w844 & w938;
assign w2073 = w827 & ~w1661;
assign w2074 = w1626 & ~w1857;
assign w2075 = (~w2071 & w2070) | (~w2071 & w9726) | (w2070 & w9726);
assign w2076 = ~w2072 & ~w2073;
assign w2077 = ~w2074 & w2076;
assign w2078 = w2075 & w2077;
assign w2079 = pi1108 & w863;
assign w2080 = pi1068 & w861;
assign w2081 = pi1735 & w865;
assign w2082 = pi1014 & w859;
assign w2083 = ~w2079 & ~w2080;
assign w2084 = ~w2081 & ~w2082;
assign w2085 = w2083 & w2084;
assign w2086 = ~pi0316 & w870;
assign w2087 = w934 & ~w1974;
assign w2088 = pi1004 & w865;
assign w2089 = pi1665 & w859;
assign w2090 = pi1628 & w861;
assign w2091 = pi1258 & w863;
assign w2092 = ~w2088 & ~w2089;
assign w2093 = ~w2090 & ~w2091;
assign w2094 = w2092 & w2093;
assign w2095 = w1838 & ~w2094;
assign w2096 = w873 & ~w2011;
assign w2097 = (~w2086 & w2085) | (~w2086 & w9727) | (w2085 & w9727);
assign w2098 = ~w2087 & ~w2095;
assign w2099 = ~w2096 & w2098;
assign w2100 = w2097 & w2099;
assign w2101 = ~pi0317 & w824;
assign w2102 = w812 & ~w1624;
assign w2103 = w938 & ~w1997;
assign w2104 = pi1737 & w819;
assign w2105 = pi1296 & w813;
assign w2106 = pi1385 & w817;
assign w2107 = pi1651 & w815;
assign w2108 = ~w2104 & ~w2105;
assign w2109 = ~w2106 & ~w2107;
assign w2110 = w2108 & w2109;
assign w2111 = w1626 & ~w2110;
assign w2112 = (~w2101 & w1616) | (~w2101 & w9728) | (w1616 & w9728);
assign w2113 = ~w2102 & ~w2103;
assign w2114 = ~w2111 & w2113;
assign w2115 = w2112 & w2114;
assign w2116 = ~pi0318 & w870;
assign w2117 = w873 & ~w1953;
assign w2118 = w934 & ~w1887;
assign w2119 = pi1254 & w863;
assign w2120 = pi1661 & w859;
assign w2121 = pi1624 & w861;
assign w2122 = pi1814 & w865;
assign w2123 = ~w2119 & ~w2120;
assign w2124 = ~w2121 & ~w2122;
assign w2125 = w2123 & w2124;
assign w2126 = w1838 & ~w2125;
assign w2127 = (~w2116 & w2049) | (~w2116 & w9729) | (w2049 & w9729);
assign w2128 = ~w2117 & ~w2118;
assign w2129 = ~w2126 & w2128;
assign w2130 = w2127 & w2129;
assign w2131 = ~pi0319 & w824;
assign w2132 = w827 & ~w2070;
assign w2133 = ~w852 & w938;
assign w2134 = w812 & ~w844;
assign w2135 = (~w2131 & w1777) | (~w2131 & w9730) | (w1777 & w9730);
assign w2136 = ~w2132 & ~w2133;
assign w2137 = ~w2134 & w2136;
assign w2138 = w2135 & w2137;
assign w2139 = pi1650 & w859;
assign w2140 = pi1736 & w865;
assign w2141 = pi1616 & w861;
assign w2142 = pi1242 & w863;
assign w2143 = ~w2139 & ~w2140;
assign w2144 = ~w2141 & ~w2142;
assign w2145 = w2143 & w2144;
assign w2146 = ~pi0320 & w870;
assign w2147 = w934 & ~w2049;
assign w2148 = pi1783 & w865;
assign w2149 = pi1629 & w861;
assign w2150 = pi1666 & w859;
assign w2151 = pi1259 & w863;
assign w2152 = ~w2148 & ~w2149;
assign w2153 = ~w2150 & ~w2151;
assign w2154 = w2152 & w2153;
assign w2155 = w1838 & ~w2154;
assign w2156 = w873 & ~w2041;
assign w2157 = (~w2146 & w2145) | (~w2146 & w9731) | (w2145 & w9731);
assign w2158 = ~w2147 & ~w2155;
assign w2159 = ~w2156 & w2158;
assign w2160 = w2157 & w2159;
assign w2161 = ~pi0321 & w824;
assign w2162 = w827 & ~w1653;
assign w2163 = w938 & ~w2070;
assign w2164 = pi1000 & w819;
assign w2165 = pi1653 & w815;
assign w2166 = pi1272 & w817;
assign w2167 = pi1297 & w813;
assign w2168 = ~w2164 & ~w2165;
assign w2169 = ~w2166 & ~w2167;
assign w2170 = w2168 & w2169;
assign w2171 = w1626 & ~w2170;
assign w2172 = (~w2161 & w1661) | (~w2161 & w9732) | (w1661 & w9732);
assign w2173 = ~w2162 & ~w2163;
assign w2174 = ~w2171 & w2173;
assign w2175 = w2172 & w2174;
assign w2176 = pi1224 & w859;
assign w2177 = pi1631 & w861;
assign w2178 = pi1006 & w865;
assign w2179 = pi1261 & w863;
assign w2180 = ~w2176 & ~w2177;
assign w2181 = ~w2178 & ~w2179;
assign w2182 = w2180 & w2181;
assign w2183 = ~pi0322 & w870;
assign w2184 = w1838 & ~w2011;
assign w2185 = ~w880 & w934;
assign w2186 = ~w869 & w873;
assign w2187 = (~w2183 & w2182) | (~w2183 & w9733) | (w2182 & w9733);
assign w2188 = ~w2184 & ~w2185;
assign w2189 = ~w2186 & w2188;
assign w2190 = w2187 & w2189;
assign w2191 = pi1007 & w865;
assign w2192 = pi1263 & w863;
assign w2193 = pi1226 & w859;
assign w2194 = pi1633 & w861;
assign w2195 = ~w2191 & ~w2192;
assign w2196 = ~w2193 & ~w2194;
assign w2197 = w2195 & w2196;
assign w2198 = ~pi0323 & w870;
assign w2199 = ~w898 & w934;
assign w2200 = w1838 & ~w2041;
assign w2201 = w873 & ~w890;
assign w2202 = (~w2198 & w2197) | (~w2198 & w9734) | (w2197 & w9734);
assign w2203 = ~w2199 & ~w2200;
assign w2204 = ~w2201 & w2203;
assign w2205 = w2202 & w2204;
assign w2206 = ~pi0324 & w870;
assign w2207 = w1838 & ~w2085;
assign w2208 = w873 & ~w2182;
assign w2209 = w858 & ~w1820;
assign w2210 = (~w2206 & w869) | (~w2206 & w9735) | (w869 & w9735);
assign w2211 = ~w2207 & ~w2208;
assign w2212 = ~w2209 & w2211;
assign w2213 = w2210 & w2212;
assign w2214 = ~pi0325 & w870;
assign w2215 = w1838 & ~w2145;
assign w2216 = w873 & ~w2197;
assign w2217 = w858 & ~w1895;
assign w2218 = (~w2214 & w890) | (~w2214 & w9736) | (w890 & w9736);
assign w2219 = ~w2215 & ~w2216;
assign w2220 = ~w2217 & w2219;
assign w2221 = w2218 & w2220;
assign w2222 = ~pi0326 & w870;
assign w2223 = w934 & ~w2182;
assign w2224 = w858 & ~w1836;
assign w2225 = pi1026 & w859;
assign w2226 = pi1618 & w861;
assign w2227 = pi1246 & w863;
assign w2228 = pi1738 & w865;
assign w2229 = ~w2225 & ~w2226;
assign w2230 = ~w2227 & ~w2228;
assign w2231 = w2229 & w2230;
assign w2232 = w1838 & ~w2231;
assign w2233 = (~w2222 & w1820) | (~w2222 & w9737) | (w1820 & w9737);
assign w2234 = ~w2223 & ~w2224;
assign w2235 = ~w2232 & w2234;
assign w2236 = w2233 & w2235;
assign w2237 = ~pi0327 & w870;
assign w2238 = w934 & ~w2197;
assign w2239 = w873 & ~w1895;
assign w2240 = pi1049 & w861;
assign w2241 = pi1247 & w863;
assign w2242 = pi1739 & w865;
assign w2243 = pi1654 & w859;
assign w2244 = ~w2240 & ~w2241;
assign w2245 = ~w2242 & ~w2243;
assign w2246 = w2244 & w2245;
assign w2247 = w1838 & ~w2246;
assign w2248 = (~w2237 & w1879) | (~w2237 & w9738) | (w1879 & w9738);
assign w2249 = ~w2238 & ~w2239;
assign w2250 = ~w2247 & w2249;
assign w2251 = w2248 & w2250;
assign w2252 = pi0812 & pi2032;
assign w2253 = ~pi0322 & ~pi2032;
assign w2254 = ~w2252 & ~w2253;
assign w2255 = ~pi2247 & w522;
assign w2256 = ~pi2249 & w532;
assign w2257 = ~pi1155 & ~pi2008;
assign w2258 = pi1155 & pi2008;
assign w2259 = ~pi1154 & ~pi2137;
assign w2260 = ~w2258 & w2259;
assign w2261 = ~pi2020 & ~w2257;
assign w2262 = ~w2260 & w2261;
assign w2263 = pi1150 & ~w2262;
assign w2264 = ~w2262 & w9739;
assign w2265 = (~pi0332 & w2262) | (~pi0332 & w9741) | (w2262 & w9741);
assign w2266 = ~pi2254 & ~w2265;
assign w2267 = pi0333 & pi2059;
assign w2268 = pi0840 & ~pi2059;
assign w2269 = ~w2267 & ~w2268;
assign w2270 = pi0334 & pi2057;
assign w2271 = pi0840 & ~pi2057;
assign w2272 = ~w2270 & ~w2271;
assign w2273 = pi0335 & pi2058;
assign w2274 = pi0840 & ~pi2058;
assign w2275 = ~w2273 & ~w2274;
assign w2276 = pi0336 & pi2056;
assign w2277 = pi0840 & ~pi2056;
assign w2278 = ~w2276 & ~w2277;
assign w2279 = w602 & w9742;
assign w2280 = ~pi1020 & pi1165;
assign w2281 = w2279 & w2280;
assign w2282 = pi0214 & pi0236;
assign w2283 = pi1369 & w2282;
assign w2284 = ~pi0214 & ~pi0236;
assign w2285 = pi1673 & w2284;
assign w2286 = ~pi0214 & pi0236;
assign w2287 = pi1319 & w2286;
assign w2288 = pi0214 & ~pi0236;
assign w2289 = pi1344 & w2288;
assign w2290 = ~w2283 & ~w2285;
assign w2291 = ~w2287 & ~w2289;
assign w2292 = w2290 & w2291;
assign w2293 = (pi1035 & ~w602) | (pi1035 & w9743) | (~w602 & w9743);
assign w2294 = ~pi0337 & w2293;
assign w2295 = pi1020 & ~pi1165;
assign w2296 = w2279 & w2295;
assign w2297 = pi1355 & w2288;
assign w2298 = pi1380 & w2282;
assign w2299 = pi1330 & w2286;
assign w2300 = pi1681 & w2284;
assign w2301 = ~w2297 & ~w2298;
assign w2302 = ~w2299 & ~w2300;
assign w2303 = w2301 & w2302;
assign w2304 = w2296 & ~w2303;
assign w2305 = (~w2294 & w2292) | (~w2294 & w9744) | (w2292 & w9744);
assign w2306 = ~w2304 & w2305;
assign w2307 = w613 & w9745;
assign w2308 = pi1171 & ~pi1789;
assign w2309 = w2307 & w2308;
assign w2310 = pi0215 & ~pi0238;
assign w2311 = pi1419 & w2310;
assign w2312 = pi1395 & w610;
assign w2313 = ~pi0215 & ~pi0238;
assign w2314 = pi1688 & w2313;
assign w2315 = pi1444 & w714;
assign w2316 = ~w2311 & ~w2312;
assign w2317 = ~w2314 & ~w2315;
assign w2318 = w2316 & w2317;
assign w2319 = (pi1169 & ~w613) | (pi1169 & w9746) | (~w613 & w9746);
assign w2320 = ~pi0338 & w2319;
assign w2321 = ~pi1171 & pi1789;
assign w2322 = w2307 & w2321;
assign w2323 = pi1406 & w610;
assign w2324 = pi1696 & w2313;
assign w2325 = pi1430 & w2310;
assign w2326 = pi1456 & w714;
assign w2327 = ~w2323 & ~w2324;
assign w2328 = ~w2325 & ~w2326;
assign w2329 = w2327 & w2328;
assign w2330 = w2322 & ~w2329;
assign w2331 = (~w2320 & w2318) | (~w2320 & w9747) | (w2318 & w9747);
assign w2332 = ~w2330 & w2331;
assign w2333 = pi1386 & w610;
assign w2334 = pi1796 & w2313;
assign w2335 = pi1436 & w714;
assign w2336 = pi1411 & w2310;
assign w2337 = ~w2333 & ~w2334;
assign w2338 = ~w2335 & ~w2336;
assign w2339 = w2337 & w2338;
assign w2340 = ~pi0339 & w2319;
assign w2341 = pi1811 & w714;
assign w2342 = pi1822 & w610;
assign w2343 = pi1694 & w2313;
assign w2344 = pi1817 & w2310;
assign w2345 = ~w2341 & ~w2342;
assign w2346 = ~w2343 & ~w2344;
assign w2347 = w2345 & w2346;
assign w2348 = w2322 & ~w2347;
assign w2349 = (~w2340 & w2339) | (~w2340 & w9748) | (w2339 & w9748);
assign w2350 = ~w2348 & w2349;
assign w2351 = pi1335 & w2288;
assign w2352 = pi1668 & w2284;
assign w2353 = pi1360 & w2282;
assign w2354 = pi1310 & w2286;
assign w2355 = ~w2351 & ~w2352;
assign w2356 = ~w2353 & ~w2354;
assign w2357 = w2355 & w2356;
assign w2358 = ~pi0340 & w2293;
assign w2359 = pi1378 & w2282;
assign w2360 = pi1353 & w2288;
assign w2361 = pi1679 & w2284;
assign w2362 = pi1328 & w2286;
assign w2363 = ~w2359 & ~w2360;
assign w2364 = ~w2361 & ~w2362;
assign w2365 = w2363 & w2364;
assign w2366 = w2296 & ~w2365;
assign w2367 = (~w2358 & w2357) | (~w2358 & w9749) | (w2357 & w9749);
assign w2368 = ~w2366 & w2367;
assign w2369 = ~pi2246 & w545;
assign w2370 = ~pi2248 & w555;
assign w2371 = ~pi2250 & w565;
assign w2372 = ~pi2251 & w575;
assign w2373 = w605 & w2279;
assign w2374 = ~pi0345 & w2293;
assign w2375 = pi1356 & w2288;
assign w2376 = pi1381 & w2282;
assign w2377 = pi0959 & w2284;
assign w2378 = pi1331 & w2286;
assign w2379 = ~w2375 & ~w2376;
assign w2380 = ~w2377 & ~w2378;
assign w2381 = w2379 & w2380;
assign w2382 = w2296 & ~w2381;
assign w2383 = pi0353 & pi1035;
assign w2384 = w603 & w9750;
assign w2385 = pi0954 & w2284;
assign w2386 = pi1040 & w2282;
assign w2387 = pi1018 & w2288;
assign w2388 = pi1061 & w2286;
assign w2389 = ~w2385 & ~w2386;
assign w2390 = ~w2387 & ~w2388;
assign w2391 = w2389 & w2390;
assign w2392 = w2384 & ~w2391;
assign w2393 = w2281 & ~w2365;
assign w2394 = (~w2374 & w2357) | (~w2374 & w9751) | (w2357 & w9751);
assign w2395 = ~w2382 & ~w2392;
assign w2396 = ~w2393 & w2395;
assign w2397 = w2394 & w2396;
assign w2398 = ~pi1138 & ~pi1152;
assign w2399 = ~pi0635 & w2398;
assign w2400 = pi0929 & pi1943;
assign w2401 = ~pi1834 & w2400;
assign w2402 = ~w2399 & w2401;
assign w2403 = w2402 & w9752;
assign w2404 = w2402 & w9754;
assign w2405 = (w2402 & w9755) | (w2402 & w9756) | (w9755 & w9756);
assign w2406 = ~w2404 & w2405;
assign w2407 = ~pi1160 & ~pi2017;
assign w2408 = pi1160 & pi2017;
assign w2409 = ~pi1159 & ~pi2136;
assign w2410 = ~w2408 & w2409;
assign w2411 = ~pi2033 & ~w2407;
assign w2412 = ~w2410 & w2411;
assign w2413 = pi1145 & ~w2412;
assign w2414 = ~w2412 & w9757;
assign w2415 = (~pi0347 & w2412) | (~pi0347 & w9759) | (w2412 & w9759);
assign w2416 = ~pi2252 & ~w2415;
assign w2417 = ~pi1148 & ~pi2016;
assign w2418 = pi1148 & pi2016;
assign w2419 = ~pi1147 & ~pi2135;
assign w2420 = ~w2418 & w2419;
assign w2421 = ~pi2055 & ~w2417;
assign w2422 = ~w2420 & w2421;
assign w2423 = pi1036 & ~w2422;
assign w2424 = ~w2422 & w9760;
assign w2425 = (~pi0348 & w2422) | (~pi0348 & w9762) | (w2422 & w9762);
assign w2426 = ~pi2253 & ~w2425;
assign w2427 = ~pi0349 & w2319;
assign w2428 = w2322 & ~w2339;
assign w2429 = ~w2427 & ~w2428;
assign w2430 = ~pi0350 & w2319;
assign w2431 = ~w2318 & w2322;
assign w2432 = ~w2430 & ~w2431;
assign w2433 = ~pi0351 & w2293;
assign w2434 = ~w2292 & w2296;
assign w2435 = ~w2433 & ~w2434;
assign w2436 = ~pi0352 & w2293;
assign w2437 = w2296 & ~w2357;
assign w2438 = ~w2436 & ~w2437;
assign w2439 = (w2383 & ~w603) | (w2383 & w9763) | (~w603 & w9763);
assign w2440 = ~w2373 & ~w2439;
assign w2441 = w612 & w2307;
assign w2442 = pi0354 & pi1169;
assign w2443 = (w2442 & ~w614) | (w2442 & w9764) | (~w614 & w9764);
assign w2444 = ~w2441 & ~w2443;
assign w2445 = w2402 & w9765;
assign w2446 = pi1138 & ~pi1152;
assign w2447 = pi0197 & w2446;
assign w2448 = pi1901 & w2398;
assign w2449 = ~w2447 & ~w2448;
assign w2450 = w2445 & ~w2449;
assign w2451 = (~pi0355 & ~w2402) | (~pi0355 & w9766) | (~w2402 & w9766);
assign w2452 = ~w2450 & ~w2451;
assign w2453 = pi0193 & w2446;
assign w2454 = pi1875 & w2398;
assign w2455 = ~w2453 & ~w2454;
assign w2456 = w2445 & ~w2455;
assign w2457 = (~pi0356 & ~w2402) | (~pi0356 & w9767) | (~w2402 & w9767);
assign w2458 = ~w2456 & ~w2457;
assign w2459 = w2402 & w9768;
assign w2460 = ~w2449 & w2459;
assign w2461 = (~pi0357 & ~w2402) | (~pi0357 & w9769) | (~w2402 & w9769);
assign w2462 = ~w2460 & ~w2461;
assign w2463 = ~w2455 & w2459;
assign w2464 = (~pi0358 & ~w2402) | (~pi0358 & w9770) | (~w2402 & w9770);
assign w2465 = ~w2463 & ~w2464;
assign w2466 = w2402 & w9772;
assign w2467 = (~pi0359 & ~w2402) | (~pi0359 & w9773) | (~w2402 & w9773);
assign w2468 = ~w2466 & ~w2467;
assign w2469 = w2402 & w9774;
assign w2470 = (~pi0360 & ~w2402) | (~pi0360 & w9775) | (~w2402 & w9775);
assign w2471 = ~w2469 & ~w2470;
assign w2472 = w2402 & w9776;
assign w2473 = (~pi0361 & ~w2402) | (~pi0361 & w9777) | (~w2402 & w9777);
assign w2474 = ~w2472 & ~w2473;
assign w2475 = w2402 & w9778;
assign w2476 = (~pi0362 & ~w2402) | (~pi0362 & w9779) | (~w2402 & w9779);
assign w2477 = ~w2475 & ~w2476;
assign w2478 = w2402 & w9780;
assign w2479 = (~pi0363 & ~w2402) | (~pi0363 & w9781) | (~w2402 & w9781);
assign w2480 = ~w2478 & ~w2479;
assign w2481 = w2402 & w9782;
assign w2482 = (~pi0364 & ~w2402) | (~pi0364 & w9783) | (~w2402 & w9783);
assign w2483 = ~w2481 & ~w2482;
assign w2484 = w2402 & w9784;
assign w2485 = (~pi0365 & ~w2402) | (~pi0365 & w9785) | (~w2402 & w9785);
assign w2486 = ~w2484 & ~w2485;
assign w2487 = w2402 & w9786;
assign w2488 = (~pi0366 & ~w2402) | (~pi0366 & w9787) | (~w2402 & w9787);
assign w2489 = ~w2487 & ~w2488;
assign w2490 = w2402 & w9788;
assign w2491 = (~pi0367 & ~w2402) | (~pi0367 & w9789) | (~w2402 & w9789);
assign w2492 = ~w2490 & ~w2491;
assign w2493 = w2402 & w9790;
assign w2494 = (~pi0368 & ~w2402) | (~pi0368 & w9791) | (~w2402 & w9791);
assign w2495 = ~w2493 & ~w2494;
assign w2496 = w2402 & w9792;
assign w2497 = (~pi0369 & ~w2402) | (~pi0369 & w9793) | (~w2402 & w9793);
assign w2498 = ~w2496 & ~w2497;
assign w2499 = w2402 & w9794;
assign w2500 = ~pi0370 & ~w2459;
assign w2501 = ~w2499 & ~w2500;
assign w2502 = w2402 & w9795;
assign w2503 = ~w2449 & w2502;
assign w2504 = (~pi0371 & ~w2402) | (~pi0371 & w9796) | (~w2402 & w9796);
assign w2505 = ~w2503 & ~w2504;
assign w2506 = ~w2455 & w2502;
assign w2507 = (~pi0372 & ~w2402) | (~pi0372 & w9797) | (~w2402 & w9797);
assign w2508 = ~w2506 & ~w2507;
assign w2509 = w2402 & w9799;
assign w2510 = (~pi0373 & ~w2402) | (~pi0373 & w9800) | (~w2402 & w9800);
assign w2511 = ~w2509 & ~w2510;
assign w2512 = w2402 & w9801;
assign w2513 = (~pi0374 & ~w2402) | (~pi0374 & w9802) | (~w2402 & w9802);
assign w2514 = ~w2512 & ~w2513;
assign w2515 = w2402 & w9803;
assign w2516 = (~pi0375 & ~w2402) | (~pi0375 & w9804) | (~w2402 & w9804);
assign w2517 = ~w2515 & ~w2516;
assign w2518 = w2402 & w9805;
assign w2519 = (~pi0376 & ~w2402) | (~pi0376 & w9806) | (~w2402 & w9806);
assign w2520 = ~w2518 & ~w2519;
assign w2521 = w2402 & w9807;
assign w2522 = (~pi0377 & ~w2402) | (~pi0377 & w9808) | (~w2402 & w9808);
assign w2523 = ~w2521 & ~w2522;
assign w2524 = w2402 & w9809;
assign w2525 = (~pi0378 & ~w2402) | (~pi0378 & w9810) | (~w2402 & w9810);
assign w2526 = ~w2524 & ~w2525;
assign w2527 = w2402 & w9811;
assign w2528 = (~pi0379 & ~w2402) | (~pi0379 & w9812) | (~w2402 & w9812);
assign w2529 = ~w2527 & ~w2528;
assign w2530 = w2402 & w9813;
assign w2531 = (~pi0380 & ~w2402) | (~pi0380 & w9814) | (~w2402 & w9814);
assign w2532 = ~w2530 & ~w2531;
assign w2533 = w2402 & w9815;
assign w2534 = (~pi0381 & ~w2402) | (~pi0381 & w9816) | (~w2402 & w9816);
assign w2535 = ~w2533 & ~w2534;
assign w2536 = w2402 & w9817;
assign w2537 = (~pi0382 & ~w2402) | (~pi0382 & w9818) | (~w2402 & w9818);
assign w2538 = ~w2536 & ~w2537;
assign w2539 = w2402 & w9819;
assign w2540 = (~pi0383 & ~w2402) | (~pi0383 & w9820) | (~w2402 & w9820);
assign w2541 = ~w2539 & ~w2540;
assign w2542 = w2402 & w9821;
assign w2543 = ~pi0384 & ~w2502;
assign w2544 = ~w2542 & ~w2543;
assign w2545 = w2403 & ~w2449;
assign w2546 = (~pi0385 & ~w2402) | (~pi0385 & w9822) | (~w2402 & w9822);
assign w2547 = ~w2545 & ~w2546;
assign w2548 = w2403 & ~w2455;
assign w2549 = (~pi0386 & ~w2402) | (~pi0386 & w9823) | (~w2402 & w9823);
assign w2550 = ~w2548 & ~w2549;
assign w2551 = w2402 & w9825;
assign w2552 = (~pi0387 & ~w2402) | (~pi0387 & w9826) | (~w2402 & w9826);
assign w2553 = ~w2551 & ~w2552;
assign w2554 = w2402 & w9827;
assign w2555 = (~pi0388 & ~w2402) | (~pi0388 & w9828) | (~w2402 & w9828);
assign w2556 = ~w2554 & ~w2555;
assign w2557 = w2402 & w9829;
assign w2558 = (~pi0389 & ~w2402) | (~pi0389 & w9830) | (~w2402 & w9830);
assign w2559 = ~w2557 & ~w2558;
assign w2560 = w2402 & w9831;
assign w2561 = (~pi0390 & ~w2402) | (~pi0390 & w9832) | (~w2402 & w9832);
assign w2562 = ~w2560 & ~w2561;
assign w2563 = w2402 & w9833;
assign w2564 = (~pi0391 & ~w2402) | (~pi0391 & w9834) | (~w2402 & w9834);
assign w2565 = ~w2563 & ~w2564;
assign w2566 = w2402 & w9835;
assign w2567 = (~pi0392 & ~w2402) | (~pi0392 & w9836) | (~w2402 & w9836);
assign w2568 = ~w2566 & ~w2567;
assign w2569 = w2402 & w9837;
assign w2570 = (~pi0393 & ~w2402) | (~pi0393 & w9838) | (~w2402 & w9838);
assign w2571 = ~w2569 & ~w2570;
assign w2572 = w2402 & w9839;
assign w2573 = (~pi0394 & ~w2402) | (~pi0394 & w9840) | (~w2402 & w9840);
assign w2574 = ~w2572 & ~w2573;
assign w2575 = w2402 & w9841;
assign w2576 = (~pi0395 & ~w2402) | (~pi0395 & w9842) | (~w2402 & w9842);
assign w2577 = ~w2575 & ~w2576;
assign w2578 = w2402 & w9843;
assign w2579 = (~pi0396 & ~w2402) | (~pi0396 & w9844) | (~w2402 & w9844);
assign w2580 = ~w2578 & ~w2579;
assign w2581 = w2402 & w9845;
assign w2582 = (~pi0397 & ~w2402) | (~pi0397 & w9846) | (~w2402 & w9846);
assign w2583 = ~w2581 & ~w2582;
assign w2584 = w2402 & w9847;
assign w2585 = ~pi0398 & ~w2403;
assign w2586 = ~w2584 & ~w2585;
assign w2587 = pi1875 & w2446;
assign w2588 = ~pi1138 & pi1152;
assign w2589 = pi0923 & w2588;
assign w2590 = pi0803 & w2398;
assign w2591 = ~w2587 & ~w2589;
assign w2592 = ~w2590 & w2591;
assign w2593 = w2403 & ~w2592;
assign w2594 = (~pi0399 & ~w2402) | (~pi0399 & w9848) | (~w2402 & w9848);
assign w2595 = ~w2593 & ~w2594;
assign w2596 = pi0794 & w2398;
assign w2597 = pi0814 & w2446;
assign w2598 = pi0335 & w2588;
assign w2599 = ~w2596 & ~w2597;
assign w2600 = ~w2598 & w2599;
assign w2601 = w2459 & ~w2600;
assign w2602 = (~pi0400 & ~w2402) | (~pi0400 & w9849) | (~w2402 & w9849);
assign w2603 = ~w2601 & ~w2602;
assign w2604 = pi0480 & w2446;
assign w2605 = pi0233 & w2588;
assign w2606 = pi0795 & w2398;
assign w2607 = ~w2604 & ~w2605;
assign w2608 = ~w2606 & w2607;
assign w2609 = w2459 & ~w2608;
assign w2610 = (~pi0401 & ~w2402) | (~pi0401 & w9850) | (~w2402 & w9850);
assign w2611 = ~w2609 & ~w2610;
assign w2612 = pi1935 & w2398;
assign w2613 = pi0213 & w2446;
assign w2614 = pi0197 & w2588;
assign w2615 = ~w2612 & ~w2613;
assign w2616 = ~w2614 & w2615;
assign w2617 = w2459 & ~w2616;
assign w2618 = (~pi0402 & ~w2402) | (~pi0402 & w9851) | (~w2402 & w9851);
assign w2619 = ~w2617 & ~w2618;
assign w2620 = pi0208 & w2446;
assign w2621 = pi0193 & w2588;
assign w2622 = pi1926 & w2398;
assign w2623 = ~w2620 & ~w2621;
assign w2624 = ~w2622 & w2623;
assign w2625 = w2502 & ~w2624;
assign w2626 = (~pi0403 & ~w2402) | (~pi0403 & w9852) | (~w2402 & w9852);
assign w2627 = ~w2625 & ~w2626;
assign w2628 = pi0798 & w2398;
assign w2629 = pi1961 & w2446;
assign w2630 = pi1978 & w2588;
assign w2631 = ~w2628 & ~w2629;
assign w2632 = ~w2630 & w2631;
assign w2633 = w2502 & ~w2632;
assign w2634 = (~pi0404 & ~w2402) | (~pi0404 & w9853) | (~w2402 & w9853);
assign w2635 = ~w2633 & ~w2634;
assign w2636 = w2502 & ~w2592;
assign w2637 = (~pi0405 & ~w2402) | (~pi0405 & w9854) | (~w2402 & w9854);
assign w2638 = ~w2636 & ~w2637;
assign w2639 = pi0657 & w2398;
assign w2640 = pi0947 & w2446;
assign w2641 = pi0877 & w2588;
assign w2642 = ~w2639 & ~w2640;
assign w2643 = ~w2641 & w2642;
assign w2644 = w2502 & ~w2643;
assign w2645 = (~pi0406 & ~w2402) | (~pi0406 & w9855) | (~w2402 & w9855);
assign w2646 = ~w2644 & ~w2645;
assign w2647 = w2403 & ~w2616;
assign w2648 = (~pi0407 & ~w2402) | (~pi0407 & w9856) | (~w2402 & w9856);
assign w2649 = ~w2647 & ~w2648;
assign w2650 = w2403 & ~w2624;
assign w2651 = (~pi0408 & ~w2402) | (~pi0408 & w9857) | (~w2402 & w9857);
assign w2652 = ~w2650 & ~w2651;
assign w2653 = pi1926 & w2446;
assign w2654 = pi1875 & w2588;
assign w2655 = pi0801 & w2398;
assign w2656 = ~w2653 & ~w2654;
assign w2657 = ~w2655 & w2656;
assign w2658 = w2403 & ~w2657;
assign w2659 = (~pi0409 & ~w2402) | (~pi0409 & w9858) | (~w2402 & w9858);
assign w2660 = ~w2658 & ~w2659;
assign w2661 = pi1901 & w2446;
assign w2662 = pi0947 & w2588;
assign w2663 = pi0802 & w2398;
assign w2664 = ~w2661 & ~w2662;
assign w2665 = ~w2663 & w2664;
assign w2666 = w2403 & ~w2665;
assign w2667 = (~pi0410 & ~w2402) | (~pi0410 & w9859) | (~w2402 & w9859);
assign w2668 = ~w2666 & ~w2667;
assign w2669 = ~pi0411 & ~w2402;
assign w2670 = (pi1150 & ~w2402) | (pi1150 & w9860) | (~w2402 & w9860);
assign w2671 = ~w2669 & w2670;
assign w2672 = (~pi0412 & ~w2402) | (~pi0412 & w9765) | (~w2402 & w9765);
assign w2673 = pi1150 & ~w2403;
assign w2674 = ~w2672 & w2673;
assign w2675 = pi1669 & w2284;
assign w2676 = pi1311 & w2286;
assign w2677 = pi1336 & w2288;
assign w2678 = pi1361 & w2282;
assign w2679 = ~w2675 & ~w2676;
assign w2680 = ~w2677 & ~w2678;
assign w2681 = w2679 & w2680;
assign w2682 = ~pi0413 & w2293;
assign w2683 = pi1359 & w2288;
assign w2684 = pi1384 & w2282;
assign w2685 = pi1334 & w2286;
assign w2686 = pi1683 & w2284;
assign w2687 = ~w2683 & ~w2684;
assign w2688 = ~w2685 & ~w2686;
assign w2689 = w2687 & w2688;
assign w2690 = w2281 & ~w2689;
assign w2691 = pi1382 & w2282;
assign w2692 = pi1792 & w2284;
assign w2693 = pi1357 & w2288;
assign w2694 = pi1332 & w2286;
assign w2695 = ~w2691 & ~w2692;
assign w2696 = ~w2693 & ~w2694;
assign w2697 = w2695 & w2696;
assign w2698 = w2373 & ~w2697;
assign w2699 = pi0956 & w2284;
assign w2700 = pi1372 & w2282;
assign w2701 = pi1322 & w2286;
assign w2702 = pi1347 & w2288;
assign w2703 = ~w2699 & ~w2700;
assign w2704 = ~w2701 & ~w2702;
assign w2705 = w2703 & w2704;
assign w2706 = w2384 & ~w2705;
assign w2707 = (~w2682 & w2681) | (~w2682 & w9861) | (w2681 & w9861);
assign w2708 = ~w2690 & ~w2698;
assign w2709 = ~w2706 & w2708;
assign w2710 = w2707 & w2709;
assign w2711 = pi1670 & w2284;
assign w2712 = pi1337 & w2288;
assign w2713 = pi1362 & w2282;
assign w2714 = pi1312 & w2286;
assign w2715 = ~w2711 & ~w2712;
assign w2716 = ~w2713 & ~w2714;
assign w2717 = w2715 & w2716;
assign w2718 = ~pi0414 & w2293;
assign w2719 = pi1338 & w2288;
assign w2720 = pi0952 & w2284;
assign w2721 = pi1363 & w2282;
assign w2722 = pi1313 & w2286;
assign w2723 = ~w2719 & ~w2720;
assign w2724 = ~w2721 & ~w2722;
assign w2725 = w2723 & w2724;
assign w2726 = w2296 & ~w2725;
assign w2727 = pi0961 & w2284;
assign w2728 = pi1054 & w2286;
assign w2729 = pi1039 & w2288;
assign w2730 = pi1027 & w2282;
assign w2731 = ~w2727 & ~w2728;
assign w2732 = ~w2729 & ~w2730;
assign w2733 = w2731 & w2732;
assign w2734 = w2373 & ~w2733;
assign w2735 = pi1374 & w2282;
assign w2736 = pi1324 & w2286;
assign w2737 = pi1675 & w2284;
assign w2738 = pi1349 & w2288;
assign w2739 = ~w2735 & ~w2736;
assign w2740 = ~w2737 & ~w2738;
assign w2741 = w2739 & w2740;
assign w2742 = w2384 & ~w2741;
assign w2743 = (~w2718 & w2717) | (~w2718 & w9862) | (w2717 & w9862);
assign w2744 = ~w2726 & ~w2734;
assign w2745 = ~w2742 & w2744;
assign w2746 = w2743 & w2745;
assign w2747 = pi1314 & w2286;
assign w2748 = pi0953 & w2284;
assign w2749 = pi1364 & w2282;
assign w2750 = pi1339 & w2288;
assign w2751 = ~w2747 & ~w2748;
assign w2752 = ~w2749 & ~w2750;
assign w2753 = w2751 & w2752;
assign w2754 = ~pi0415 & w2293;
assign w2755 = pi1065 & w2286;
assign w2756 = pi1052 & w2288;
assign w2757 = pi1041 & w2282;
assign w2758 = pi1818 & w2284;
assign w2759 = ~w2755 & ~w2756;
assign w2760 = ~w2757 & ~w2758;
assign w2761 = w2759 & w2760;
assign w2762 = w2281 & ~w2761;
assign w2763 = w2373 & ~w2681;
assign w2764 = pi1678 & w2284;
assign w2765 = pi1325 & w2286;
assign w2766 = pi1375 & w2282;
assign w2767 = pi1350 & w2288;
assign w2768 = ~w2764 & ~w2765;
assign w2769 = ~w2766 & ~w2767;
assign w2770 = w2768 & w2769;
assign w2771 = w2384 & ~w2770;
assign w2772 = (~w2754 & w2753) | (~w2754 & w9863) | (w2753 & w9863);
assign w2773 = ~w2762 & ~w2763;
assign w2774 = ~w2771 & w2773;
assign w2775 = w2772 & w2774;
assign w2776 = pi1365 & w2282;
assign w2777 = pi1340 & w2288;
assign w2778 = pi1671 & w2284;
assign w2779 = pi1315 & w2286;
assign w2780 = ~w2776 & ~w2777;
assign w2781 = ~w2778 & ~w2779;
assign w2782 = w2780 & w2781;
assign w2783 = ~pi0416 & w2293;
assign w2784 = w2281 & ~w2725;
assign w2785 = w2373 & ~w2717;
assign w2786 = pi1056 & w2286;
assign w2787 = pi1033 & w2282;
assign w2788 = pi1045 & w2288;
assign w2789 = pi1676 & w2284;
assign w2790 = ~w2786 & ~w2787;
assign w2791 = ~w2788 & ~w2789;
assign w2792 = w2790 & w2791;
assign w2793 = w2384 & ~w2792;
assign w2794 = (~w2783 & w2782) | (~w2783 & w9864) | (w2782 & w9864);
assign w2795 = ~w2784 & ~w2785;
assign w2796 = ~w2793 & w2795;
assign w2797 = w2794 & w2796;
assign w2798 = ~pi0417 & w2293;
assign w2799 = w2296 & ~w2391;
assign w2800 = w2373 & ~w2761;
assign w2801 = pi1677 & w2284;
assign w2802 = pi1326 & w2286;
assign w2803 = pi1376 & w2282;
assign w2804 = pi1351 & w2288;
assign w2805 = ~w2801 & ~w2802;
assign w2806 = ~w2803 & ~w2804;
assign w2807 = w2805 & w2806;
assign w2808 = w2384 & ~w2807;
assign w2809 = (~w2798 & w2753) | (~w2798 & w9865) | (w2753 & w9865);
assign w2810 = ~w2799 & ~w2800;
assign w2811 = ~w2808 & w2810;
assign w2812 = w2809 & w2811;
assign w2813 = ~pi0418 & w2293;
assign w2814 = w2281 & ~w2733;
assign w2815 = pi0960 & w2284;
assign w2816 = pi1383 & w2282;
assign w2817 = pi1333 & w2286;
assign w2818 = pi1358 & w2288;
assign w2819 = ~w2815 & ~w2816;
assign w2820 = ~w2817 & ~w2818;
assign w2821 = w2819 & w2820;
assign w2822 = w2373 & ~w2821;
assign w2823 = pi1060 & w2286;
assign w2824 = pi1032 & w2282;
assign w2825 = pi1046 & w2288;
assign w2826 = pi1806 & w2284;
assign w2827 = ~w2823 & ~w2824;
assign w2828 = ~w2825 & ~w2826;
assign w2829 = w2827 & w2828;
assign w2830 = w2384 & ~w2829;
assign w2831 = (~w2813 & w2717) | (~w2813 & w9866) | (w2717 & w9866);
assign w2832 = ~w2814 & ~w2822;
assign w2833 = ~w2830 & w2832;
assign w2834 = w2831 & w2833;
assign w2835 = pi1672 & w2284;
assign w2836 = pi1342 & w2288;
assign w2837 = pi1317 & w2286;
assign w2838 = pi1367 & w2282;
assign w2839 = ~w2835 & ~w2836;
assign w2840 = ~w2837 & ~w2838;
assign w2841 = w2839 & w2840;
assign w2842 = ~pi0419 & w2293;
assign w2843 = w2373 & ~w2753;
assign w2844 = pi1053 & w2286;
assign w2845 = pi1029 & w2282;
assign w2846 = pi1799 & w2284;
assign w2847 = pi1044 & w2288;
assign w2848 = ~w2844 & ~w2845;
assign w2849 = ~w2846 & ~w2847;
assign w2850 = w2848 & w2849;
assign w2851 = w2384 & ~w2850;
assign w2852 = w2281 & ~w2391;
assign w2853 = (~w2842 & w2841) | (~w2842 & w9867) | (w2841 & w9867);
assign w2854 = ~w2843 & ~w2851;
assign w2855 = ~w2852 & w2854;
assign w2856 = w2853 & w2855;
assign w2857 = ~pi0420 & w2293;
assign w2858 = w2281 & ~w2681;
assign w2859 = w2373 & ~w2689;
assign w2860 = pi0957 & w2284;
assign w2861 = pi1373 & w2282;
assign w2862 = pi1323 & w2286;
assign w2863 = pi1348 & w2288;
assign w2864 = ~w2860 & ~w2861;
assign w2865 = ~w2862 & ~w2863;
assign w2866 = w2864 & w2865;
assign w2867 = w2384 & ~w2866;
assign w2868 = (~w2857 & w2761) | (~w2857 & w9868) | (w2761 & w9868);
assign w2869 = ~w2858 & ~w2859;
assign w2870 = ~w2867 & w2869;
assign w2871 = w2868 & w2870;
assign w2872 = pi0955 & w2284;
assign w2873 = pi1368 & w2282;
assign w2874 = pi1318 & w2286;
assign w2875 = pi1343 & w2288;
assign w2876 = ~w2872 & ~w2873;
assign w2877 = ~w2874 & ~w2875;
assign w2878 = w2876 & w2877;
assign w2879 = ~pi0421 & w2293;
assign w2880 = pi1316 & w2286;
assign w2881 = pi1808 & w2284;
assign w2882 = pi1341 & w2288;
assign w2883 = pi1366 & w2282;
assign w2884 = ~w2880 & ~w2881;
assign w2885 = ~w2882 & ~w2883;
assign w2886 = w2884 & w2885;
assign w2887 = w2281 & ~w2886;
assign w2888 = pi0958 & w2284;
assign w2889 = pi1354 & w2288;
assign w2890 = pi1329 & w2286;
assign w2891 = pi1379 & w2282;
assign w2892 = ~w2888 & ~w2889;
assign w2893 = ~w2890 & ~w2891;
assign w2894 = w2892 & w2893;
assign w2895 = w2384 & ~w2894;
assign w2896 = w2373 & ~w2782;
assign w2897 = (~w2879 & w2878) | (~w2879 & w9869) | (w2878 & w9869);
assign w2898 = ~w2887 & ~w2895;
assign w2899 = ~w2896 & w2898;
assign w2900 = w2897 & w2899;
assign w2901 = ~pi0422 & w2293;
assign w2902 = w2296 & ~w2886;
assign w2903 = w2373 & ~w2725;
assign w2904 = pi1327 & w2286;
assign w2905 = pi1680 & w2284;
assign w2906 = pi1352 & w2288;
assign w2907 = pi1377 & w2282;
assign w2908 = ~w2904 & ~w2905;
assign w2909 = ~w2906 & ~w2907;
assign w2910 = w2908 & w2909;
assign w2911 = w2384 & ~w2910;
assign w2912 = (~w2901 & w2782) | (~w2901 & w9870) | (w2782 & w9870);
assign w2913 = ~w2902 & ~w2903;
assign w2914 = ~w2911 & w2913;
assign w2915 = w2912 & w2914;
assign w2916 = ~pi0423 & w2293;
assign w2917 = pi1042 & w2288;
assign w2918 = pi1055 & w2286;
assign w2919 = pi1682 & w2284;
assign w2920 = pi1028 & w2282;
assign w2921 = ~w2917 & ~w2918;
assign w2922 = ~w2919 & ~w2920;
assign w2923 = w2921 & w2922;
assign w2924 = w2296 & ~w2923;
assign w2925 = ~w2292 & w2373;
assign w2926 = w2281 & ~w2303;
assign w2927 = (~w2916 & w2886) | (~w2916 & w9871) | (w2886 & w9871);
assign w2928 = ~w2924 & ~w2925;
assign w2929 = ~w2926 & w2928;
assign w2930 = w2927 & w2929;
assign w2931 = ~pi0424 & w2293;
assign w2932 = ~w2365 & w2373;
assign w2933 = w2296 & ~w2697;
assign w2934 = w2384 & ~w2841;
assign w2935 = (~w2931 & w2381) | (~w2931 & w9872) | (w2381 & w9872);
assign w2936 = ~w2932 & ~w2933;
assign w2937 = ~w2934 & w2936;
assign w2938 = w2935 & w2937;
assign w2939 = ~pi0425 & w2293;
assign w2940 = ~w2303 & w2373;
assign w2941 = w2296 & ~w2821;
assign w2942 = w2384 & ~w2878;
assign w2943 = (~w2939 & w2923) | (~w2939 & w9873) | (w2923 & w9873);
assign w2944 = ~w2940 & ~w2941;
assign w2945 = ~w2942 & w2944;
assign w2946 = w2943 & w2945;
assign w2947 = ~pi0426 & w2293;
assign w2948 = w2296 & ~w2689;
assign w2949 = w2373 & ~w2381;
assign w2950 = pi1370 & w2282;
assign w2951 = pi1320 & w2286;
assign w2952 = pi1345 & w2288;
assign w2953 = pi1815 & w2284;
assign w2954 = ~w2950 & ~w2951;
assign w2955 = ~w2952 & ~w2953;
assign w2956 = w2954 & w2955;
assign w2957 = w2384 & ~w2956;
assign w2958 = (~w2947 & w2697) | (~w2947 & w9874) | (w2697 & w9874);
assign w2959 = ~w2948 & ~w2949;
assign w2960 = ~w2957 & w2959;
assign w2961 = w2958 & w2960;
assign w2962 = ~pi0427 & w2293;
assign w2963 = w2296 & ~w2733;
assign w2964 = w2373 & ~w2923;
assign w2965 = pi1321 & w2286;
assign w2966 = pi1674 & w2284;
assign w2967 = pi1346 & w2288;
assign w2968 = pi1371 & w2282;
assign w2969 = ~w2965 & ~w2966;
assign w2970 = ~w2967 & ~w2968;
assign w2971 = w2969 & w2970;
assign w2972 = w2384 & ~w2971;
assign w2973 = (~w2962 & w2821) | (~w2962 & w9875) | (w2821 & w9875);
assign w2974 = ~w2963 & ~w2964;
assign w2975 = ~w2972 & w2974;
assign w2976 = w2973 & w2975;
assign w2977 = pi1408 & w610;
assign w2978 = pi1433 & w2310;
assign w2979 = pi1766 & w2313;
assign w2980 = pi1458 & w714;
assign w2981 = ~w2977 & ~w2978;
assign w2982 = ~w2979 & ~w2980;
assign w2983 = w2981 & w2982;
assign w2984 = ~pi0428 & w2319;
assign w2985 = pi1412 & w2310;
assign w2986 = pi1437 & w714;
assign w2987 = pi1387 & w610;
assign w2988 = pi1684 & w2313;
assign w2989 = ~w2985 & ~w2986;
assign w2990 = ~w2987 & ~w2988;
assign w2991 = w2989 & w2990;
assign w2992 = w2322 & ~w2991;
assign w2993 = pi1698 & w2313;
assign w2994 = pi1829 & w610;
assign w2995 = pi1805 & w2310;
assign w2996 = pi1801 & w714;
assign w2997 = ~w2993 & ~w2994;
assign w2998 = ~w2995 & ~w2996;
assign w2999 = w2997 & w2998;
assign w3000 = w2309 & ~w2999;
assign w3001 = w614 & w9876;
assign w3002 = pi0966 & w2313;
assign w3003 = pi1021 & w610;
assign w3004 = pi1826 & w2310;
assign w3005 = pi1812 & w714;
assign w3006 = ~w3002 & ~w3003;
assign w3007 = ~w3004 & ~w3005;
assign w3008 = w3006 & w3007;
assign w3009 = w3001 & ~w3008;
assign w3010 = (~w2984 & w2983) | (~w2984 & w9877) | (w2983 & w9877);
assign w3011 = ~w2992 & ~w3000;
assign w3012 = ~w3009 & w3011;
assign w3013 = w3010 & w3012;
assign w3014 = pi1460 & w714;
assign w3015 = pi1435 & w2310;
assign w3016 = pi0971 & w2313;
assign w3017 = pi1410 & w610;
assign w3018 = ~w3014 & ~w3015;
assign w3019 = ~w3016 & ~w3017;
assign w3020 = w3018 & w3019;
assign w3021 = ~pi0429 & w2319;
assign w3022 = pi1434 & w2310;
assign w3023 = pi0970 & w2313;
assign w3024 = pi1409 & w610;
assign w3025 = pi1459 & w714;
assign w3026 = ~w3022 & ~w3023;
assign w3027 = ~w3024 & ~w3025;
assign w3028 = w3026 & w3027;
assign w3029 = w2441 & ~w3028;
assign w3030 = pi1823 & w2310;
assign w3031 = pi1685 & w2313;
assign w3032 = pi1024 & w610;
assign w3033 = pi1816 & w714;
assign w3034 = ~w3030 & ~w3031;
assign w3035 = ~w3032 & ~w3033;
assign w3036 = w3034 & w3035;
assign w3037 = w2322 & ~w3036;
assign w3038 = pi1422 & w2310;
assign w3039 = pi1770 & w2313;
assign w3040 = pi1448 & w714;
assign w3041 = pi1398 & w610;
assign w3042 = ~w3038 & ~w3039;
assign w3043 = ~w3040 & ~w3041;
assign w3044 = w3042 & w3043;
assign w3045 = w3001 & ~w3044;
assign w3046 = (~w3021 & w3020) | (~w3021 & w9878) | (w3020 & w9878);
assign w3047 = ~w3029 & ~w3037;
assign w3048 = ~w3045 & w3047;
assign w3049 = w3046 & w3048;
assign w3050 = ~pi0430 & w2319;
assign w3051 = w2309 & ~w2991;
assign w3052 = pi1388 & w610;
assign w3053 = pi1413 & w2310;
assign w3054 = pi1790 & w2313;
assign w3055 = pi1438 & w714;
assign w3056 = ~w3052 & ~w3053;
assign w3057 = ~w3054 & ~w3055;
assign w3058 = w3056 & w3057;
assign w3059 = w2322 & ~w3058;
assign w3060 = pi1449 & w714;
assign w3061 = pi1399 & w610;
assign w3062 = pi0967 & w2313;
assign w3063 = pi1423 & w2310;
assign w3064 = ~w3060 & ~w3061;
assign w3065 = ~w3062 & ~w3063;
assign w3066 = w3064 & w3065;
assign w3067 = w3001 & ~w3066;
assign w3068 = (~w3050 & w2999) | (~w3050 & w9879) | (w2999 & w9879);
assign w3069 = ~w3051 & ~w3059;
assign w3070 = ~w3067 & w3069;
assign w3071 = w3068 & w3070;
assign w3072 = pi1440 & w714;
assign w3073 = pi1415 & w2310;
assign w3074 = pi0963 & w2313;
assign w3075 = pi1390 & w610;
assign w3076 = ~w3072 & ~w3073;
assign w3077 = ~w3074 & ~w3075;
assign w3078 = w3076 & w3077;
assign w3079 = ~pi0431 & w2319;
assign w3080 = w2441 & ~w2991;
assign w3081 = w2309 & ~w3058;
assign w3082 = pi1019 & w610;
assign w3083 = pi1810 & w714;
assign w3084 = pi1691 & w2313;
assign w3085 = pi1819 & w2310;
assign w3086 = ~w3082 & ~w3083;
assign w3087 = ~w3084 & ~w3085;
assign w3088 = w3086 & w3087;
assign w3089 = w3001 & ~w3088;
assign w3090 = (~w3079 & w3078) | (~w3079 & w9880) | (w3078 & w9880);
assign w3091 = ~w3080 & ~w3081;
assign w3092 = ~w3089 & w3091;
assign w3093 = w3090 & w3092;
assign w3094 = ~pi0432 & w2319;
assign w3095 = pi1827 & w2310;
assign w3096 = pi1813 & w714;
assign w3097 = pi1022 & w610;
assign w3098 = pi1686 & w2313;
assign w3099 = ~w3095 & ~w3096;
assign w3100 = ~w3097 & ~w3098;
assign w3101 = w3099 & w3100;
assign w3102 = w2322 & ~w3101;
assign w3103 = pi1414 & w2310;
assign w3104 = pi0962 & w2313;
assign w3105 = pi1439 & w714;
assign w3106 = pi1389 & w610;
assign w3107 = ~w3103 & ~w3104;
assign w3108 = ~w3105 & ~w3106;
assign w3109 = w3107 & w3108;
assign w3110 = w2309 & ~w3109;
assign w3111 = pi1401 & w610;
assign w3112 = pi1425 & w2310;
assign w3113 = pi1451 & w714;
assign w3114 = pi1692 & w2313;
assign w3115 = ~w3111 & ~w3112;
assign w3116 = ~w3113 & ~w3114;
assign w3117 = w3115 & w3116;
assign w3118 = w3001 & ~w3117;
assign w3119 = (~w3094 & w3036) | (~w3094 & w9881) | (w3036 & w9881);
assign w3120 = ~w3102 & ~w3110;
assign w3121 = ~w3118 & w3120;
assign w3122 = w3119 & w3121;
assign w3123 = pi1441 & w714;
assign w3124 = pi0964 & w2313;
assign w3125 = pi1392 & w610;
assign w3126 = pi1416 & w2310;
assign w3127 = ~w3123 & ~w3124;
assign w3128 = ~w3125 & ~w3126;
assign w3129 = w3127 & w3128;
assign w3130 = ~pi0433 & w2319;
assign w3131 = w2441 & ~w3058;
assign w3132 = w2309 & ~w3078;
assign w3133 = pi1402 & w610;
assign w3134 = pi1426 & w2310;
assign w3135 = pi1778 & w2313;
assign w3136 = pi1452 & w714;
assign w3137 = ~w3133 & ~w3134;
assign w3138 = ~w3135 & ~w3136;
assign w3139 = w3137 & w3138;
assign w3140 = w3001 & ~w3139;
assign w3141 = (~w3130 & w3129) | (~w3130 & w9882) | (w3129 & w9882);
assign w3142 = ~w3131 & ~w3132;
assign w3143 = ~w3140 & w3142;
assign w3144 = w3141 & w3143;
assign w3145 = pi1687 & w2313;
assign w3146 = pi1443 & w714;
assign w3147 = pi1394 & w610;
assign w3148 = pi1418 & w2310;
assign w3149 = ~w3145 & ~w3146;
assign w3150 = ~w3147 & ~w3148;
assign w3151 = w3149 & w3150;
assign w3152 = ~pi0434 & w2319;
assign w3153 = w2309 & ~w3129;
assign w3154 = pi1769 & w2313;
assign w3155 = pi1428 & w2310;
assign w3156 = pi1454 & w714;
assign w3157 = pi1404 & w610;
assign w3158 = ~w3154 & ~w3155;
assign w3159 = ~w3156 & ~w3157;
assign w3160 = w3158 & w3159;
assign w3161 = w3001 & ~w3160;
assign w3162 = w2441 & ~w3078;
assign w3163 = (~w3152 & w3151) | (~w3152 & w9883) | (w3151 & w9883);
assign w3164 = ~w3153 & ~w3161;
assign w3165 = ~w3162 & w3164;
assign w3166 = w3163 & w3165;
assign w3167 = pi1809 & w714;
assign w3168 = pi1023 & w610;
assign w3169 = pi1825 & w2310;
assign w3170 = pi0965 & w2313;
assign w3171 = ~w3167 & ~w3168;
assign w3172 = ~w3169 & ~w3170;
assign w3173 = w3171 & w3172;
assign w3174 = ~pi0435 & w2319;
assign w3175 = w2441 & ~w3101;
assign w3176 = pi1455 & w714;
assign w3177 = pi1405 & w610;
assign w3178 = pi1429 & w2310;
assign w3179 = pi0968 & w2313;
assign w3180 = ~w3176 & ~w3177;
assign w3181 = ~w3178 & ~w3179;
assign w3182 = w3180 & w3181;
assign w3183 = w3001 & ~w3182;
assign w3184 = pi1442 & w714;
assign w3185 = pi1393 & w610;
assign w3186 = pi1417 & w2310;
assign w3187 = pi1788 & w2313;
assign w3188 = ~w3184 & ~w3185;
assign w3189 = ~w3186 & ~w3187;
assign w3190 = w3188 & w3189;
assign w3191 = w2309 & ~w3190;
assign w3192 = (~w3174 & w3173) | (~w3174 & w9884) | (w3173 & w9884);
assign w3193 = ~w3175 & ~w3183;
assign w3194 = ~w3191 & w3193;
assign w3195 = w3192 & w3194;
assign w3196 = pi0969 & w2313;
assign w3197 = pi1803 & w714;
assign w3198 = pi1830 & w610;
assign w3199 = pi1431 & w2310;
assign w3200 = ~w3196 & ~w3197;
assign w3201 = ~w3198 & ~w3199;
assign w3202 = w3200 & w3201;
assign w3203 = ~pi0436 & w2319;
assign w3204 = ~w2339 & w2441;
assign w3205 = w3001 & ~w3129;
assign w3206 = w2309 & ~w2347;
assign w3207 = (~w3203 & w3202) | (~w3203 & w9885) | (w3202 & w9885);
assign w3208 = ~w3204 & ~w3205;
assign w3209 = ~w3206 & w3208;
assign w3210 = w3207 & w3209;
assign w3211 = ~pi0437 & w2319;
assign w3212 = pi1432 & w2310;
assign w3213 = pi1407 & w610;
assign w3214 = pi1457 & w714;
assign w3215 = pi1697 & w2313;
assign w3216 = ~w3212 & ~w3213;
assign w3217 = ~w3214 & ~w3215;
assign w3218 = w3216 & w3217;
assign w3219 = w2322 & ~w3218;
assign w3220 = ~w2318 & w2441;
assign w3221 = w2309 & ~w2329;
assign w3222 = (~w3211 & w3190) | (~w3211 & w9886) | (w3190 & w9886);
assign w3223 = ~w3219 & ~w3220;
assign w3224 = ~w3221 & w3223;
assign w3225 = w3222 & w3224;
assign w3226 = ~pi0438 & w2319;
assign w3227 = w3001 & ~w3151;
assign w3228 = w2309 & ~w3202;
assign w3229 = w2322 & ~w2983;
assign w3230 = (~w3226 & w2347) | (~w3226 & w9887) | (w2347 & w9887);
assign w3231 = ~w3227 & ~w3228;
assign w3232 = ~w3229 & w3231;
assign w3233 = w3230 & w3232;
assign w3234 = ~pi0439 & w2319;
assign w3235 = w2322 & ~w2999;
assign w3236 = w2441 & ~w3202;
assign w3237 = pi1782 & w2313;
assign w3238 = pi1445 & w714;
assign w3239 = pi1420 & w2310;
assign w3240 = pi1396 & w610;
assign w3241 = ~w3237 & ~w3238;
assign w3242 = ~w3239 & ~w3240;
assign w3243 = w3241 & w3242;
assign w3244 = w3001 & ~w3243;
assign w3245 = (~w3234 & w2983) | (~w3234 & w9888) | (w2983 & w9888);
assign w3246 = ~w3235 & ~w3236;
assign w3247 = ~w3244 & w3246;
assign w3248 = w3245 & w3247;
assign w3249 = ~pi0440 & w2319;
assign w3250 = w2441 & ~w3218;
assign w3251 = w2309 & ~w3028;
assign w3252 = pi1446 & w714;
assign w3253 = pi1689 & w2313;
assign w3254 = pi1421 & w2310;
assign w3255 = pi1397 & w610;
assign w3256 = ~w3252 & ~w3253;
assign w3257 = ~w3254 & ~w3255;
assign w3258 = w3256 & w3257;
assign w3259 = w3001 & ~w3258;
assign w3260 = (~w3249 & w3020) | (~w3249 & w9889) | (w3020 & w9889);
assign w3261 = ~w3250 & ~w3251;
assign w3262 = ~w3259 & w3261;
assign w3263 = w3260 & w3262;
assign w3264 = pi1979 & w2446;
assign w3265 = pi1962 & w2588;
assign w3266 = pi0791 & w2398;
assign w3267 = ~w3264 & ~w3265;
assign w3268 = ~w3266 & w3267;
assign w3269 = w2445 & ~w3268;
assign w3270 = (~pi0441 & ~w2402) | (~pi0441 & w9890) | (~w2402 & w9890);
assign w3271 = ~w3269 & ~w3270;
assign w3272 = pi0814 & w2588;
assign w3273 = pi0877 & w2446;
assign w3274 = pi0792 & w2398;
assign w3275 = ~w3272 & ~w3273;
assign w3276 = ~w3274 & w3275;
assign w3277 = w2445 & ~w3276;
assign w3278 = (~pi0442 & ~w2402) | (~pi0442 & w9891) | (~w2402 & w9891);
assign w3279 = ~w3277 & ~w3278;
assign w3280 = pi0871 & w2446;
assign w3281 = pi0480 & w2588;
assign w3282 = pi0793 & w2398;
assign w3283 = ~w3280 & ~w3281;
assign w3284 = ~w3282 & w3283;
assign w3285 = w2445 & ~w3284;
assign w3286 = (~pi0443 & ~w2402) | (~pi0443 & w9892) | (~w2402 & w9892);
assign w3287 = ~w3285 & ~w3286;
assign w3288 = w2445 & ~w2600;
assign w3289 = (~pi0444 & ~w2402) | (~pi0444 & w9893) | (~w2402 & w9893);
assign w3290 = ~w3288 & ~w3289;
assign w3291 = w2445 & ~w2608;
assign w3292 = (~pi0445 & ~w2402) | (~pi0445 & w9894) | (~w2402 & w9894);
assign w3293 = ~w3291 & ~w3292;
assign w3294 = pi0335 & w2446;
assign w3295 = pi0213 & w2588;
assign w3296 = pi0796 & w2398;
assign w3297 = ~w3294 & ~w3295;
assign w3298 = ~w3296 & w3297;
assign w3299 = w2445 & ~w3298;
assign w3300 = (~pi0446 & ~w2402) | (~pi0446 & w9895) | (~w2402 & w9895);
assign w3301 = ~w3299 & ~w3300;
assign w3302 = pi0233 & w2446;
assign w3303 = pi0208 & w2588;
assign w3304 = pi0797 & w2398;
assign w3305 = ~w3302 & ~w3303;
assign w3306 = ~w3304 & w3305;
assign w3307 = w2445 & ~w3306;
assign w3308 = (~pi0447 & ~w2402) | (~pi0447 & w9896) | (~w2402 & w9896);
assign w3309 = ~w3307 & ~w3308;
assign w3310 = w2445 & ~w2632;
assign w3311 = (~pi0448 & ~w2402) | (~pi0448 & w9897) | (~w2402 & w9897);
assign w3312 = ~w3310 & ~w3311;
assign w3313 = pi1144 & pi1905;
assign w3314 = ~pi0946 & pi1930;
assign w3315 = (pi0449 & ~w3314) | (pi0449 & w9898) | (~w3314 & w9898);
assign w3316 = ~w3313 & ~w3315;
assign w3317 = w629 & w9899;
assign w3318 = pi0450 & ~w3317;
assign w3319 = w637 & w9900;
assign w3320 = pi0451 & ~w3319;
assign w3321 = w645 & w9901;
assign w3322 = pi0452 & ~w3321;
assign w3323 = w621 & w9902;
assign w3324 = pi0453 & ~w3323;
assign w3325 = ~pi0454 & w2319;
assign w3326 = w2309 & ~w3218;
assign w3327 = w3001 & ~w3173;
assign w3328 = ~w2329 & w2441;
assign w3329 = (~w3325 & w3028) | (~w3325 & w9903) | (w3028 & w9903);
assign w3330 = ~w3326 & ~w3327;
assign w3331 = ~w3328 & w3330;
assign w3332 = w3329 & w3331;
assign w3333 = ~pi0455 & w2319;
assign w3334 = w2322 & ~w3190;
assign w3335 = w2309 & ~w3101;
assign w3336 = pi1453 & w714;
assign w3337 = pi1695 & w2313;
assign w3338 = pi1427 & w2310;
assign w3339 = pi1403 & w610;
assign w3340 = ~w3336 & ~w3337;
assign w3341 = ~w3338 & ~w3339;
assign w3342 = w3340 & w3341;
assign w3343 = w3001 & ~w3342;
assign w3344 = (~w3333 & w3109) | (~w3333 & w9904) | (w3109 & w9904);
assign w3345 = ~w3334 & ~w3335;
assign w3346 = ~w3343 & w3345;
assign w3347 = w3344 & w3346;
assign w3348 = ~pi0457 & w2319;
assign w3349 = w2322 & ~w3109;
assign w3350 = w2441 & ~w3020;
assign w3351 = pi1400 & w610;
assign w3352 = pi1450 & w714;
assign w3353 = pi1424 & w2310;
assign w3354 = pi1693 & w2313;
assign w3355 = ~w3351 & ~w3352;
assign w3356 = ~w3353 & ~w3354;
assign w3357 = w3355 & w3356;
assign w3358 = w3001 & ~w3357;
assign w3359 = (~w3348 & w3036) | (~w3348 & w9905) | (w3036 & w9905);
assign w3360 = ~w3349 & ~w3350;
assign w3361 = ~w3358 & w3360;
assign w3362 = w3359 & w3361;
assign w3363 = ~pi1134 & ~pi1146;
assign w3364 = ~pi0790 & w3363;
assign w3365 = pi0939 & pi1952;
assign w3366 = ~pi1876 & w3365;
assign w3367 = ~w3364 & w3366;
assign w3368 = w3367 & w9906;
assign w3369 = pi1134 & ~pi1146;
assign w3370 = pi0196 & w3369;
assign w3371 = pi1886 & w3363;
assign w3372 = ~w3370 & ~w3371;
assign w3373 = w3368 & ~w3372;
assign w3374 = (~pi0458 & ~w3367) | (~pi0458 & w9907) | (~w3367 & w9907);
assign w3375 = ~w3373 & ~w3374;
assign w3376 = w3367 & w9908;
assign w3377 = w3367 & w9910;
assign w3378 = (~pi0459 & ~w3367) | (~pi0459 & w9911) | (~w3367 & w9911);
assign w3379 = ~w3377 & ~w3378;
assign w3380 = w3367 & w9912;
assign w3381 = (~pi0460 & ~w3367) | (~pi0460 & w9913) | (~w3367 & w9913);
assign w3382 = ~w3380 & ~w3381;
assign w3383 = ~pi1157 & ~pi1158;
assign w3384 = ~pi0821 & w3383;
assign w3385 = pi0938 & ~pi1931;
assign w3386 = pi1881 & w3385;
assign w3387 = ~w3384 & w3386;
assign w3388 = w3387 & w9914;
assign w3389 = w3387 & w9916;
assign w3390 = (~pi0461 & ~w3387) | (~pi0461 & w9917) | (~w3387 & w9917);
assign w3391 = ~w3389 & ~w3390;
assign w3392 = w3387 & w9918;
assign w3393 = (~pi0462 & ~w3387) | (~pi0462 & w9919) | (~w3387 & w9919);
assign w3394 = ~w3392 & ~w3393;
assign w3395 = w3367 & w9921;
assign w3396 = (w3367 & w9922) | (w3367 & w9923) | (w9922 & w9923);
assign w3397 = ~w3395 & w3396;
assign w3398 = w3387 & w9924;
assign w3399 = (~pi0464 & ~w3387) | (~pi0464 & w9925) | (~w3387 & w9925);
assign w3400 = ~w3398 & ~w3399;
assign w3401 = w3387 & w9926;
assign w3402 = w3387 & w9928;
assign w3403 = (~pi0465 & ~w3387) | (~pi0465 & w9929) | (~w3387 & w9929);
assign w3404 = ~w3402 & ~w3403;
assign w3405 = w3387 & w9930;
assign w3406 = (~pi0466 & ~w3387) | (~pi0466 & w9931) | (~w3387 & w9931);
assign w3407 = ~w3405 & ~w3406;
assign w3408 = w3387 & w9932;
assign w3409 = (~pi0467 & ~w3387) | (~pi0467 & w9933) | (~w3387 & w9933);
assign w3410 = ~w3408 & ~w3409;
assign w3411 = w3387 & w9934;
assign w3412 = w3387 & w9936;
assign w3413 = (~pi0468 & ~w3387) | (~pi0468 & w9937) | (~w3387 & w9937);
assign w3414 = ~w3412 & ~w3413;
assign w3415 = w3387 & w9938;
assign w3416 = (~pi0469 & ~w3387) | (~pi0469 & w9939) | (~w3387 & w9939);
assign w3417 = ~w3415 & ~w3416;
assign w3418 = w3387 & w9940;
assign w3419 = (~pi0470 & ~w3387) | (~pi0470 & w9941) | (~w3387 & w9941);
assign w3420 = ~w3418 & ~w3419;
assign w3421 = w3367 & w9942;
assign w3422 = w3421 & w9943;
assign w3423 = (~pi0471 & ~w3367) | (~pi0471 & w9944) | (~w3367 & w9944);
assign w3424 = ~w3422 & ~w3423;
assign w3425 = w2403 & ~w3298;
assign w3426 = (~pi0472 & ~w2402) | (~pi0472 & w9945) | (~w2402 & w9945);
assign w3427 = ~w3425 & ~w3426;
assign w3428 = w2403 & ~w3268;
assign w3429 = (~pi0473 & ~w2402) | (~pi0473 & w9946) | (~w2402 & w9946);
assign w3430 = ~w3428 & ~w3429;
assign w3431 = w2403 & ~w2608;
assign w3432 = (~pi0474 & ~w2402) | (~pi0474 & w9947) | (~w2402 & w9947);
assign w3433 = ~w3431 & ~w3432;
assign w3434 = w3367 & w9948;
assign w3435 = ~pi1134 & pi1146;
assign w3436 = pi1983 & w3435;
assign w3437 = pi1984 & w3369;
assign w3438 = pi0831 & w3363;
assign w3439 = ~w3436 & ~w3437;
assign w3440 = ~w3438 & w3439;
assign w3441 = w3434 & ~w3440;
assign w3442 = (~pi0475 & ~w3367) | (~pi0475 & w9949) | (~w3367 & w9949);
assign w3443 = ~w3441 & ~w3442;
assign w3444 = w2459 & ~w3306;
assign w3445 = (~pi0476 & ~w2402) | (~pi0476 & w9950) | (~w2402 & w9950);
assign w3446 = ~w3444 & ~w3445;
assign w3447 = w2459 & ~w2665;
assign w3448 = (~pi0477 & ~w2402) | (~pi0477 & w9951) | (~w2402 & w9951);
assign w3449 = ~w3447 & ~w3448;
assign w3450 = pi0478 & pi2056;
assign w3451 = pi0876 & ~pi2056;
assign w3452 = ~w3450 & ~w3451;
assign w3453 = pi0479 & pi2057;
assign w3454 = pi0876 & ~pi2057;
assign w3455 = ~w3453 & ~w3454;
assign w3456 = pi0480 & pi2058;
assign w3457 = pi0876 & ~pi2058;
assign w3458 = ~w3456 & ~w3457;
assign w3459 = pi0481 & pi2059;
assign w3460 = pi0876 & ~pi2059;
assign w3461 = ~w3459 & ~w3460;
assign w3462 = ~w3372 & w3421;
assign w3463 = (~pi0482 & ~w3367) | (~pi0482 & w9952) | (~w3367 & w9952);
assign w3464 = ~w3462 & ~w3463;
assign w3465 = pi0192 & w3369;
assign w3466 = pi1852 & w3363;
assign w3467 = ~w3465 & ~w3466;
assign w3468 = w3421 & ~w3467;
assign w3469 = (~pi0483 & ~w3367) | (~pi0483 & w9953) | (~w3367 & w9953);
assign w3470 = ~w3468 & ~w3469;
assign w3471 = w3421 & w9954;
assign w3472 = (~pi0484 & ~w3367) | (~pi0484 & w9955) | (~w3367 & w9955);
assign w3473 = ~w3471 & ~w3472;
assign w3474 = w3421 & w9956;
assign w3475 = (~pi0485 & ~w3367) | (~pi0485 & w9957) | (~w3367 & w9957);
assign w3476 = ~w3474 & ~w3475;
assign w3477 = w3421 & w9958;
assign w3478 = (~pi0486 & ~w3367) | (~pi0486 & w9959) | (~w3367 & w9959);
assign w3479 = ~w3477 & ~w3478;
assign w3480 = w3387 & w9960;
assign w3481 = ~pi1157 & pi1158;
assign w3482 = pi0195 & w3481;
assign w3483 = pi1883 & w3383;
assign w3484 = ~w3482 & ~w3483;
assign w3485 = w3480 & ~w3484;
assign w3486 = (~pi0487 & ~w3387) | (~pi0487 & w9961) | (~w3387 & w9961);
assign w3487 = ~w3485 & ~w3486;
assign w3488 = pi0191 & w3481;
assign w3489 = pi1853 & w3383;
assign w3490 = ~w3488 & ~w3489;
assign w3491 = w3480 & ~w3490;
assign w3492 = (~pi0488 & ~w3387) | (~pi0488 & w9962) | (~w3387 & w9962);
assign w3493 = ~w3491 & ~w3492;
assign w3494 = w3421 & w9963;
assign w3495 = (~pi0489 & ~w3367) | (~pi0489 & w9964) | (~w3367 & w9964);
assign w3496 = ~w3494 & ~w3495;
assign w3497 = w3421 & w9965;
assign w3498 = (~pi0490 & ~w3367) | (~pi0490 & w9966) | (~w3367 & w9966);
assign w3499 = ~w3497 & ~w3498;
assign w3500 = w3421 & w9967;
assign w3501 = (~pi0491 & ~w3367) | (~pi0491 & w9968) | (~w3367 & w9968);
assign w3502 = ~w3500 & ~w3501;
assign w3503 = w3421 & w9969;
assign w3504 = (~pi0492 & ~w3367) | (~pi0492 & w9970) | (~w3367 & w9970);
assign w3505 = ~w3503 & ~w3504;
assign w3506 = w3411 & ~w3484;
assign w3507 = (~pi0493 & ~w3387) | (~pi0493 & w9971) | (~w3387 & w9971);
assign w3508 = ~w3506 & ~w3507;
assign w3509 = w3411 & ~w3490;
assign w3510 = (~pi0494 & ~w3387) | (~pi0494 & w9972) | (~w3387 & w9972);
assign w3511 = ~w3509 & ~w3510;
assign w3512 = w3387 & w9973;
assign w3513 = (~pi0495 & ~w3387) | (~pi0495 & w9974) | (~w3387 & w9974);
assign w3514 = ~w3512 & ~w3513;
assign w3515 = w3387 & w9975;
assign w3516 = (~pi0496 & ~w3387) | (~pi0496 & w9976) | (~w3387 & w9976);
assign w3517 = ~w3515 & ~w3516;
assign w3518 = w3421 & w9977;
assign w3519 = (~pi0497 & ~w3367) | (~pi0497 & w9978) | (~w3367 & w9978);
assign w3520 = ~w3518 & ~w3519;
assign w3521 = w3387 & w9979;
assign w3522 = (~pi0498 & ~w3387) | (~pi0498 & w9980) | (~w3387 & w9980);
assign w3523 = ~w3521 & ~w3522;
assign w3524 = w3387 & w9981;
assign w3525 = (~pi0499 & ~w3387) | (~pi0499 & w9982) | (~w3387 & w9982);
assign w3526 = ~w3524 & ~w3525;
assign w3527 = w3387 & w9983;
assign w3528 = (~pi0500 & ~w3387) | (~pi0500 & w9984) | (~w3387 & w9984);
assign w3529 = ~w3527 & ~w3528;
assign w3530 = w3421 & w9985;
assign w3531 = (~pi0501 & ~w3367) | (~pi0501 & w9986) | (~w3367 & w9986);
assign w3532 = ~w3530 & ~w3531;
assign w3533 = w3387 & w9987;
assign w3534 = (~pi0502 & ~w3387) | (~pi0502 & w9988) | (~w3387 & w9988);
assign w3535 = ~w3533 & ~w3534;
assign w3536 = w3387 & w9989;
assign w3537 = (~pi0503 & ~w3387) | (~pi0503 & w9990) | (~w3387 & w9990);
assign w3538 = ~w3536 & ~w3537;
assign w3539 = w3387 & w9991;
assign w3540 = (~pi0504 & ~w3387) | (~pi0504 & w9992) | (~w3387 & w9992);
assign w3541 = ~w3539 & ~w3540;
assign w3542 = w3387 & w9993;
assign w3543 = ~pi0505 & ~w3411;
assign w3544 = ~w3542 & ~w3543;
assign w3545 = w3421 & w9994;
assign w3546 = (~pi0506 & ~w3367) | (~pi0506 & w9995) | (~w3367 & w9995);
assign w3547 = ~w3545 & ~w3546;
assign w3548 = w3401 & ~w3484;
assign w3549 = (~pi0507 & ~w3387) | (~pi0507 & w9996) | (~w3387 & w9996);
assign w3550 = ~w3548 & ~w3549;
assign w3551 = w3401 & ~w3490;
assign w3552 = (~pi0508 & ~w3387) | (~pi0508 & w9997) | (~w3387 & w9997);
assign w3553 = ~w3551 & ~w3552;
assign w3554 = w3421 & w9998;
assign w3555 = ~pi0509 & ~w3421;
assign w3556 = ~w3554 & ~w3555;
assign w3557 = w3387 & w9999;
assign w3558 = (~pi0510 & ~w3387) | (~pi0510 & w10000) | (~w3387 & w10000);
assign w3559 = ~w3557 & ~w3558;
assign w3560 = w3387 & w10001;
assign w3561 = (~pi0511 & ~w3387) | (~pi0511 & w10002) | (~w3387 & w10002);
assign w3562 = ~w3560 & ~w3561;
assign w3563 = w3387 & w10003;
assign w3564 = (~pi0512 & ~w3387) | (~pi0512 & w10004) | (~w3387 & w10004);
assign w3565 = ~w3563 & ~w3564;
assign w3566 = w3387 & w10005;
assign w3567 = (~pi0513 & ~w3387) | (~pi0513 & w10006) | (~w3387 & w10006);
assign w3568 = ~w3566 & ~w3567;
assign w3569 = w3387 & w10007;
assign w3570 = (~pi0514 & ~w3387) | (~pi0514 & w10008) | (~w3387 & w10008);
assign w3571 = ~w3569 & ~w3570;
assign w3572 = w3387 & w10009;
assign w3573 = (~pi0515 & ~w3387) | (~pi0515 & w10010) | (~w3387 & w10010);
assign w3574 = ~w3572 & ~w3573;
assign w3575 = w3387 & w10011;
assign w3576 = (~pi0516 & ~w3387) | (~pi0516 & w10012) | (~w3387 & w10012);
assign w3577 = ~w3575 & ~w3576;
assign w3578 = w3387 & w10013;
assign w3579 = (~pi0517 & ~w3387) | (~pi0517 & w10014) | (~w3387 & w10014);
assign w3580 = ~w3578 & ~w3579;
assign w3581 = w3387 & w10015;
assign w3582 = ~pi0518 & ~w3401;
assign w3583 = ~w3581 & ~w3582;
assign w3584 = w3388 & ~w3484;
assign w3585 = (~pi0519 & ~w3387) | (~pi0519 & w10016) | (~w3387 & w10016);
assign w3586 = ~w3584 & ~w3585;
assign w3587 = w3388 & ~w3490;
assign w3588 = (~pi0520 & ~w3387) | (~pi0520 & w10017) | (~w3387 & w10017);
assign w3589 = ~w3587 & ~w3588;
assign w3590 = w3387 & w10018;
assign w3591 = (~pi0521 & ~w3387) | (~pi0521 & w10019) | (~w3387 & w10019);
assign w3592 = ~w3590 & ~w3591;
assign w3593 = w3387 & w10020;
assign w3594 = (~pi0522 & ~w3387) | (~pi0522 & w10021) | (~w3387 & w10021);
assign w3595 = ~w3593 & ~w3594;
assign w3596 = w3387 & w10022;
assign w3597 = (~pi0523 & ~w3387) | (~pi0523 & w10023) | (~w3387 & w10023);
assign w3598 = ~w3596 & ~w3597;
assign w3599 = w3387 & w10024;
assign w3600 = (~pi0524 & ~w3387) | (~pi0524 & w10025) | (~w3387 & w10025);
assign w3601 = ~w3599 & ~w3600;
assign w3602 = w3387 & w10026;
assign w3603 = (~pi0525 & ~w3387) | (~pi0525 & w10027) | (~w3387 & w10027);
assign w3604 = ~w3602 & ~w3603;
assign w3605 = w3387 & w10028;
assign w3606 = (~pi0526 & ~w3387) | (~pi0526 & w10029) | (~w3387 & w10029);
assign w3607 = ~w3605 & ~w3606;
assign w3608 = w3387 & w10030;
assign w3609 = (~pi0527 & ~w3387) | (~pi0527 & w10031) | (~w3387 & w10031);
assign w3610 = ~w3608 & ~w3609;
assign w3611 = w3387 & w10032;
assign w3612 = (~pi0528 & ~w3387) | (~pi0528 & w10033) | (~w3387 & w10033);
assign w3613 = ~w3611 & ~w3612;
assign w3614 = w3387 & w10034;
assign w3615 = ~pi0529 & ~w3388;
assign w3616 = ~w3614 & ~w3615;
assign w3617 = ~w3372 & w3376;
assign w3618 = (~pi0530 & ~w3367) | (~pi0530 & w10035) | (~w3367 & w10035);
assign w3619 = ~w3617 & ~w3618;
assign w3620 = w3376 & ~w3467;
assign w3621 = (~pi0531 & ~w3367) | (~pi0531 & w10036) | (~w3367 & w10036);
assign w3622 = ~w3620 & ~w3621;
assign w3623 = w3367 & w10037;
assign w3624 = (~pi0532 & ~w3367) | (~pi0532 & w10038) | (~w3367 & w10038);
assign w3625 = ~w3623 & ~w3624;
assign w3626 = w3367 & w10039;
assign w3627 = (~pi0533 & ~w3367) | (~pi0533 & w10040) | (~w3367 & w10040);
assign w3628 = ~w3626 & ~w3627;
assign w3629 = w3367 & w10041;
assign w3630 = (~pi0534 & ~w3367) | (~pi0534 & w10042) | (~w3367 & w10042);
assign w3631 = ~w3629 & ~w3630;
assign w3632 = w3367 & w10043;
assign w3633 = (~pi0535 & ~w3367) | (~pi0535 & w10044) | (~w3367 & w10044);
assign w3634 = ~w3632 & ~w3633;
assign w3635 = w3367 & w10045;
assign w3636 = (~pi0536 & ~w3367) | (~pi0536 & w10046) | (~w3367 & w10046);
assign w3637 = ~w3635 & ~w3636;
assign w3638 = w3367 & w10047;
assign w3639 = (~pi0537 & ~w3367) | (~pi0537 & w10048) | (~w3367 & w10048);
assign w3640 = ~w3638 & ~w3639;
assign w3641 = w3367 & w10049;
assign w3642 = (~pi0538 & ~w3367) | (~pi0538 & w10050) | (~w3367 & w10050);
assign w3643 = ~w3641 & ~w3642;
assign w3644 = w3367 & w10051;
assign w3645 = (~pi0539 & ~w3367) | (~pi0539 & w10052) | (~w3367 & w10052);
assign w3646 = ~w3644 & ~w3645;
assign w3647 = w3367 & w10053;
assign w3648 = (~pi0540 & ~w3367) | (~pi0540 & w10054) | (~w3367 & w10054);
assign w3649 = ~w3647 & ~w3648;
assign w3650 = w3367 & w10055;
assign w3651 = ~pi0541 & ~w3376;
assign w3652 = ~w3650 & ~w3651;
assign w3653 = w3368 & ~w3467;
assign w3654 = (~pi0542 & ~w3367) | (~pi0542 & w10056) | (~w3367 & w10056);
assign w3655 = ~w3653 & ~w3654;
assign w3656 = ~w3372 & w3434;
assign w3657 = (~pi0543 & ~w3367) | (~pi0543 & w10057) | (~w3367 & w10057);
assign w3658 = ~w3656 & ~w3657;
assign w3659 = w3434 & ~w3467;
assign w3660 = (~pi0544 & ~w3367) | (~pi0544 & w10058) | (~w3367 & w10058);
assign w3661 = ~w3659 & ~w3660;
assign w3662 = w3367 & w10060;
assign w3663 = (~pi0545 & ~w3367) | (~pi0545 & w10061) | (~w3367 & w10061);
assign w3664 = ~w3662 & ~w3663;
assign w3665 = w3367 & w10062;
assign w3666 = (~pi0546 & ~w3367) | (~pi0546 & w10063) | (~w3367 & w10063);
assign w3667 = ~w3665 & ~w3666;
assign w3668 = w3367 & w10064;
assign w3669 = (~pi0547 & ~w3367) | (~pi0547 & w10065) | (~w3367 & w10065);
assign w3670 = ~w3668 & ~w3669;
assign w3671 = w3367 & w10066;
assign w3672 = (~pi0548 & ~w3367) | (~pi0548 & w10067) | (~w3367 & w10067);
assign w3673 = ~w3671 & ~w3672;
assign w3674 = w3367 & w10068;
assign w3675 = (~pi0549 & ~w3367) | (~pi0549 & w10069) | (~w3367 & w10069);
assign w3676 = ~w3674 & ~w3675;
assign w3677 = w3367 & w10070;
assign w3678 = (~pi0550 & ~w3367) | (~pi0550 & w10071) | (~w3367 & w10071);
assign w3679 = ~w3677 & ~w3678;
assign w3680 = w3367 & w10072;
assign w3681 = (~pi0551 & ~w3367) | (~pi0551 & w10073) | (~w3367 & w10073);
assign w3682 = ~w3680 & ~w3681;
assign w3683 = w3367 & w10074;
assign w3684 = (~pi0552 & ~w3367) | (~pi0552 & w10075) | (~w3367 & w10075);
assign w3685 = ~w3683 & ~w3684;
assign w3686 = w3367 & w10076;
assign w3687 = (~pi0553 & ~w3367) | (~pi0553 & w10077) | (~w3367 & w10077);
assign w3688 = ~w3686 & ~w3687;
assign w3689 = w3367 & w10078;
assign w3690 = (~pi0554 & ~w3367) | (~pi0554 & w10079) | (~w3367 & w10079);
assign w3691 = ~w3689 & ~w3690;
assign w3692 = w3367 & w10080;
assign w3693 = (~pi0555 & ~w3367) | (~pi0555 & w10081) | (~w3367 & w10081);
assign w3694 = ~w3692 & ~w3693;
assign w3695 = w3367 & w10082;
assign w3696 = ~pi0556 & ~w3434;
assign w3697 = ~w3695 & ~w3696;
assign w3698 = w2403 & ~w2643;
assign w3699 = (~pi0557 & ~w2402) | (~pi0557 & w10083) | (~w2402 & w10083);
assign w3700 = ~w3698 & ~w3699;
assign w3701 = pi0804 & w2398;
assign w3702 = pi0871 & w2588;
assign w3703 = pi0923 & w2446;
assign w3704 = ~w3701 & ~w3702;
assign w3705 = ~w3703 & w3704;
assign w3706 = w2403 & ~w3705;
assign w3707 = (~pi0558 & ~w2402) | (~pi0558 & w10084) | (~w2402 & w10084);
assign w3708 = ~w3706 & ~w3707;
assign w3709 = pi1980 & w3435;
assign w3710 = pi1960 & w3369;
assign w3711 = pi0824 & w3363;
assign w3712 = ~w3709 & ~w3710;
assign w3713 = ~w3711 & w3712;
assign w3714 = w3421 & ~w3713;
assign w3715 = (~pi0559 & ~w3367) | (~pi0559 & w10085) | (~w3367 & w10085);
assign w3716 = ~w3714 & ~w3715;
assign w3717 = pi0822 & w3363;
assign w3718 = pi1924 & w3369;
assign w3719 = pi1852 & w3435;
assign w3720 = ~w3717 & ~w3718;
assign w3721 = ~w3719 & w3720;
assign w3722 = w3421 & ~w3721;
assign w3723 = (~pi0560 & ~w3367) | (~pi0560 & w10086) | (~w3367 & w10086);
assign w3724 = ~w3722 & ~w3723;
assign w3725 = pi0950 & w3435;
assign w3726 = pi1886 & w3369;
assign w3727 = pi0827 & w3363;
assign w3728 = ~w3725 & ~w3726;
assign w3729 = ~w3727 & w3728;
assign w3730 = w3421 & ~w3729;
assign w3731 = (~pi0561 & ~w3367) | (~pi0561 & w10087) | (~w3367 & w10087);
assign w3732 = ~w3730 & ~w3731;
assign w3733 = pi1924 & w3435;
assign w3734 = pi1980 & w3369;
assign w3735 = pi0823 & w3363;
assign w3736 = ~w3733 & ~w3734;
assign w3737 = ~w3735 & w3736;
assign w3738 = w3376 & ~w3737;
assign w3739 = (~pi0562 & ~w3367) | (~pi0562 & w10088) | (~w3367 & w10088);
assign w3740 = ~w3738 & ~w3739;
assign w3741 = pi0829 & w3363;
assign w3742 = pi0915 & w3369;
assign w3743 = pi0866 & w3435;
assign w3744 = ~w3741 & ~w3742;
assign w3745 = ~w3743 & w3744;
assign w3746 = w3421 & ~w3745;
assign w3747 = (~pi0563 & ~w3367) | (~pi0563 & w10089) | (~w3367 & w10089);
assign w3748 = ~w3746 & ~w3747;
assign w3749 = w2459 & ~w3268;
assign w3750 = (~pi0564 & ~w2402) | (~pi0564 & w10090) | (~w2402 & w10090);
assign w3751 = ~w3749 & ~w3750;
assign w3752 = w2459 & ~w3276;
assign w3753 = (~pi0565 & ~w2402) | (~pi0565 & w10091) | (~w2402 & w10091);
assign w3754 = ~w3752 & ~w3753;
assign w3755 = w2459 & ~w3284;
assign w3756 = (~pi0566 & ~w2402) | (~pi0566 & w10092) | (~w2402 & w10092);
assign w3757 = ~w3755 & ~w3756;
assign w3758 = pi1934 & w3435;
assign w3759 = pi1983 & w3369;
assign w3760 = pi0825 & w3363;
assign w3761 = ~w3758 & ~w3759;
assign w3762 = ~w3760 & w3761;
assign w3763 = w3376 & ~w3762;
assign w3764 = (~pi0567 & ~w3367) | (~pi0567 & w10093) | (~w3367 & w10093);
assign w3765 = ~w3763 & ~w3764;
assign w3766 = w3376 & ~w3745;
assign w3767 = (~pi0568 & ~w3367) | (~pi0568 & w10094) | (~w3367 & w10094);
assign w3768 = ~w3766 & ~w3767;
assign w3769 = w2459 & ~w3298;
assign w3770 = (~pi0569 & ~w2402) | (~pi0569 & w10095) | (~w2402 & w10095);
assign w3771 = ~w3769 & ~w3770;
assign w3772 = w2459 & ~w2632;
assign w3773 = (~pi0570 & ~w2402) | (~pi0570 & w10096) | (~w2402 & w10096);
assign w3774 = ~w3772 & ~w3773;
assign w3775 = pi0799 & w2398;
assign w3776 = pi1962 & w2446;
assign w3777 = pi1935 & w2588;
assign w3778 = ~w3775 & ~w3776;
assign w3779 = ~w3777 & w3778;
assign w3780 = w2459 & ~w3779;
assign w3781 = (~pi0571 & ~w2402) | (~pi0571 & w10097) | (~w2402 & w10097);
assign w3782 = ~w3780 & ~w3781;
assign w3783 = pi1978 & w2446;
assign w3784 = pi1926 & w2588;
assign w3785 = pi0800 & w2398;
assign w3786 = ~w3783 & ~w3784;
assign w3787 = ~w3785 & w3786;
assign w3788 = w2459 & ~w3787;
assign w3789 = (~pi0572 & ~w2402) | (~pi0572 & w10098) | (~w2402 & w10098);
assign w3790 = ~w3788 & ~w3789;
assign w3791 = pi1935 & w2446;
assign w3792 = pi1901 & w2588;
assign w3793 = pi0751 & w2398;
assign w3794 = ~w3791 & ~w3792;
assign w3795 = ~w3793 & w3794;
assign w3796 = w2459 & ~w3795;
assign w3797 = (~pi0573 & ~w2402) | (~pi0573 & w10099) | (~w2402 & w10099);
assign w3798 = ~w3796 & ~w3797;
assign w3799 = w2459 & ~w2657;
assign w3800 = (~pi0574 & ~w2402) | (~pi0574 & w10100) | (~w2402 & w10100);
assign w3801 = ~w3799 & ~w3800;
assign w3802 = w2459 & ~w2592;
assign w3803 = (~pi0575 & ~w2402) | (~pi0575 & w10101) | (~w2402 & w10101);
assign w3804 = ~w3802 & ~w3803;
assign w3805 = w2459 & ~w2643;
assign w3806 = (~pi0576 & ~w2402) | (~pi0576 & w10102) | (~w2402 & w10102);
assign w3807 = ~w3805 & ~w3806;
assign w3808 = w2459 & ~w3705;
assign w3809 = (~pi0577 & ~w2402) | (~pi0577 & w10103) | (~w2402 & w10103);
assign w3810 = ~w3808 & ~w3809;
assign w3811 = w2502 & ~w3268;
assign w3812 = (~pi0578 & ~w2402) | (~pi0578 & w10104) | (~w2402 & w10104);
assign w3813 = ~w3811 & ~w3812;
assign w3814 = w2502 & ~w3276;
assign w3815 = (~pi0579 & ~w2402) | (~pi0579 & w10105) | (~w2402 & w10105);
assign w3816 = ~w3814 & ~w3815;
assign w3817 = w2502 & ~w3284;
assign w3818 = (~pi0580 & ~w2402) | (~pi0580 & w10106) | (~w2402 & w10106);
assign w3819 = ~w3817 & ~w3818;
assign w3820 = w2502 & ~w2608;
assign w3821 = (~pi0581 & ~w2402) | (~pi0581 & w10107) | (~w2402 & w10107);
assign w3822 = ~w3820 & ~w3821;
assign w3823 = w2502 & ~w3298;
assign w3824 = (~pi0582 & ~w2402) | (~pi0582 & w10108) | (~w2402 & w10108);
assign w3825 = ~w3823 & ~w3824;
assign w3826 = w2502 & ~w3306;
assign w3827 = (~pi0583 & ~w2402) | (~pi0583 & w10109) | (~w2402 & w10109);
assign w3828 = ~w3826 & ~w3827;
assign w3829 = w2502 & ~w2616;
assign w3830 = (~pi0584 & ~w2402) | (~pi0584 & w10110) | (~w2402 & w10110);
assign w3831 = ~w3829 & ~w3830;
assign w3832 = w2459 & ~w2624;
assign w3833 = (~pi0585 & ~w2402) | (~pi0585 & w10111) | (~w2402 & w10111);
assign w3834 = ~w3832 & ~w3833;
assign w3835 = w2502 & ~w2600;
assign w3836 = (~pi0586 & ~w2402) | (~pi0586 & w10112) | (~w2402 & w10112);
assign w3837 = ~w3835 & ~w3836;
assign w3838 = w2502 & ~w3779;
assign w3839 = (~pi0587 & ~w2402) | (~pi0587 & w10113) | (~w2402 & w10113);
assign w3840 = ~w3838 & ~w3839;
assign w3841 = w2502 & ~w3787;
assign w3842 = (~pi0588 & ~w2402) | (~pi0588 & w10114) | (~w2402 & w10114);
assign w3843 = ~w3841 & ~w3842;
assign w3844 = w2502 & ~w2665;
assign w3845 = (~pi0589 & ~w2402) | (~pi0589 & w10115) | (~w2402 & w10115);
assign w3846 = ~w3844 & ~w3845;
assign w3847 = w2502 & ~w3795;
assign w3848 = (~pi0590 & ~w2402) | (~pi0590 & w10116) | (~w2402 & w10116);
assign w3849 = ~w3847 & ~w3848;
assign w3850 = w2502 & ~w2657;
assign w3851 = (~pi0591 & ~w2402) | (~pi0591 & w10117) | (~w2402 & w10117);
assign w3852 = ~w3850 & ~w3851;
assign w3853 = w2502 & ~w3705;
assign w3854 = (~pi0592 & ~w2402) | (~pi0592 & w10118) | (~w2402 & w10118);
assign w3855 = ~w3853 & ~w3854;
assign w3856 = w2403 & ~w3284;
assign w3857 = (~pi0593 & ~w2402) | (~pi0593 & w10119) | (~w2402 & w10119);
assign w3858 = ~w3856 & ~w3857;
assign w3859 = w2403 & ~w2600;
assign w3860 = (~pi0594 & ~w2402) | (~pi0594 & w10120) | (~w2402 & w10120);
assign w3861 = ~w3859 & ~w3860;
assign w3862 = w2403 & ~w3306;
assign w3863 = (~pi0595 & ~w2402) | (~pi0595 & w10121) | (~w2402 & w10121);
assign w3864 = ~w3862 & ~w3863;
assign w3865 = w2403 & ~w3276;
assign w3866 = (~pi0596 & ~w2402) | (~pi0596 & w10122) | (~w2402 & w10122);
assign w3867 = ~w3865 & ~w3866;
assign w3868 = w2403 & ~w3779;
assign w3869 = (~pi0597 & ~w2402) | (~pi0597 & w10123) | (~w2402 & w10123);
assign w3870 = ~w3868 & ~w3869;
assign w3871 = w2403 & ~w3787;
assign w3872 = (~pi0598 & ~w2402) | (~pi0598 & w10124) | (~w2402 & w10124);
assign w3873 = ~w3871 & ~w3872;
assign w3874 = w2403 & ~w3795;
assign w3875 = (~pi0599 & ~w2402) | (~pi0599 & w10125) | (~w2402 & w10125);
assign w3876 = ~w3874 & ~w3875;
assign w3877 = w2403 & ~w2632;
assign w3878 = (~pi0600 & ~w2402) | (~pi0600 & w10126) | (~w2402 & w10126);
assign w3879 = ~w3877 & ~w3878;
assign w3880 = ~pi0601 & ~w3367;
assign w3881 = (pi1036 & ~w3367) | (pi1036 & w10127) | (~w3367 & w10127);
assign w3882 = ~w3880 & w3881;
assign w3883 = (~pi0602 & ~w3367) | (~pi0602 & w9906) | (~w3367 & w9906);
assign w3884 = pi1036 & ~w3376;
assign w3885 = ~w3883 & w3884;
assign w3886 = w3368 & ~w3762;
assign w3887 = (~pi0603 & ~w3367) | (~pi0603 & w10128) | (~w3367 & w10128);
assign w3888 = ~w3886 & ~w3887;
assign w3889 = w2445 & ~w2657;
assign w3890 = (~pi0604 & ~w2402) | (~pi0604 & w10129) | (~w2402 & w10129);
assign w3891 = ~w3889 & ~w3890;
assign w3892 = pi0235 & w3435;
assign w3893 = pi0479 & w3369;
assign w3894 = pi0813 & w3363;
assign w3895 = ~w3892 & ~w3893;
assign w3896 = ~w3894 & w3895;
assign w3897 = w3368 & ~w3896;
assign w3898 = (~pi0605 & ~w3367) | (~pi0605 & w10130) | (~w3367 & w10130);
assign w3899 = ~w3897 & ~w3898;
assign w3900 = pi0334 & w3435;
assign w3901 = pi0819 & w3369;
assign w3902 = pi0835 & w3363;
assign w3903 = ~w3900 & ~w3901;
assign w3904 = ~w3902 & w3903;
assign w3905 = w3368 & ~w3904;
assign w3906 = (~pi0606 & ~w3367) | (~pi0606 & w10131) | (~w3367 & w10131);
assign w3907 = ~w3905 & ~w3906;
assign w3908 = w2445 & ~w2616;
assign w3909 = (~pi0607 & ~w2402) | (~pi0607 & w10132) | (~w2402 & w10132);
assign w3910 = ~w3908 & ~w3909;
assign w3911 = w2402 & w10134;
assign w3912 = (~pi0608 & ~w2402) | (~pi0608 & w10135) | (~w2402 & w10135);
assign w3913 = ~w3911 & ~w3912;
assign w3914 = w2402 & w10136;
assign w3915 = (~pi0609 & ~w2402) | (~pi0609 & w10137) | (~w2402 & w10137);
assign w3916 = ~w3914 & ~w3915;
assign w3917 = w2402 & w10138;
assign w3918 = (~pi0610 & ~w2402) | (~pi0610 & w10139) | (~w2402 & w10139);
assign w3919 = ~w3917 & ~w3918;
assign w3920 = w2402 & w10140;
assign w3921 = (~pi0611 & ~w2402) | (~pi0611 & w10141) | (~w2402 & w10141);
assign w3922 = ~w3920 & ~w3921;
assign w3923 = w2402 & w10142;
assign w3924 = (~pi0612 & ~w2402) | (~pi0612 & w10143) | (~w2402 & w10143);
assign w3925 = ~w3923 & ~w3924;
assign w3926 = w2402 & w10144;
assign w3927 = (~pi0613 & ~w2402) | (~pi0613 & w10145) | (~w2402 & w10145);
assign w3928 = ~w3926 & ~w3927;
assign w3929 = w3367 & w10147;
assign w3930 = (~pi0614 & ~w3367) | (~pi0614 & w10148) | (~w3367 & w10148);
assign w3931 = ~w3929 & ~w3930;
assign w3932 = w2402 & w10149;
assign w3933 = (~pi0615 & ~w2402) | (~pi0615 & w10150) | (~w2402 & w10150);
assign w3934 = ~w3932 & ~w3933;
assign w3935 = w2402 & w10151;
assign w3936 = (~pi0616 & ~w2402) | (~pi0616 & w10152) | (~w2402 & w10152);
assign w3937 = ~w3935 & ~w3936;
assign w3938 = w3367 & w10153;
assign w3939 = (~pi0617 & ~w3367) | (~pi0617 & w10154) | (~w3367 & w10154);
assign w3940 = ~w3938 & ~w3939;
assign w3941 = w2402 & w10155;
assign w3942 = (~pi0618 & ~w2402) | (~pi0618 & w10156) | (~w2402 & w10156);
assign w3943 = ~w3941 & ~w3942;
assign w3944 = w2402 & w10157;
assign w3945 = (~pi0619 & ~w2402) | (~pi0619 & w10158) | (~w2402 & w10158);
assign w3946 = ~w3944 & ~w3945;
assign w3947 = w2445 & ~w3779;
assign w3948 = (~pi0620 & ~w2402) | (~pi0620 & w10159) | (~w2402 & w10159);
assign w3949 = ~w3947 & ~w3948;
assign w3950 = w2402 & w10160;
assign w3951 = (~pi0621 & ~w2402) | (~pi0621 & w10161) | (~w2402 & w10161);
assign w3952 = ~w3950 & ~w3951;
assign w3953 = w2402 & w10162;
assign w3954 = ~pi0622 & ~w2445;
assign w3955 = ~w3953 & ~w3954;
assign w3956 = w2445 & ~w3787;
assign w3957 = (~pi0623 & ~w2402) | (~pi0623 & w10163) | (~w2402 & w10163);
assign w3958 = ~w3956 & ~w3957;
assign w3959 = w3367 & w10164;
assign w3960 = (~pi0624 & ~w3367) | (~pi0624 & w10165) | (~w3367 & w10165);
assign w3961 = ~w3959 & ~w3960;
assign w3962 = w2445 & ~w3795;
assign w3963 = (~pi0625 & ~w2402) | (~pi0625 & w10166) | (~w2402 & w10166);
assign w3964 = ~w3962 & ~w3963;
assign w3965 = w3367 & w10167;
assign w3966 = (~pi0626 & ~w3367) | (~pi0626 & w10168) | (~w3367 & w10168);
assign w3967 = ~w3965 & ~w3966;
assign w3968 = w3367 & w10169;
assign w3969 = (~pi0627 & ~w3367) | (~pi0627 & w10170) | (~w3367 & w10170);
assign w3970 = ~w3968 & ~w3969;
assign w3971 = w2445 & ~w2665;
assign w3972 = (~pi0628 & ~w2402) | (~pi0628 & w10171) | (~w2402 & w10171);
assign w3973 = ~w3971 & ~w3972;
assign w3974 = w3367 & w10172;
assign w3975 = (~pi0629 & ~w3367) | (~pi0629 & w10173) | (~w3367 & w10173);
assign w3976 = ~w3974 & ~w3975;
assign w3977 = w2445 & ~w2592;
assign w3978 = (~pi0630 & ~w2402) | (~pi0630 & w10174) | (~w2402 & w10174);
assign w3979 = ~w3977 & ~w3978;
assign w3980 = w2445 & ~w2643;
assign w3981 = (~pi0631 & ~w2402) | (~pi0631 & w10175) | (~w2402 & w10175);
assign w3982 = ~w3980 & ~w3981;
assign w3983 = w3367 & w10176;
assign w3984 = (~pi0632 & ~w3367) | (~pi0632 & w10177) | (~w3367 & w10177);
assign w3985 = ~w3983 & ~w3984;
assign w3986 = w2445 & ~w3705;
assign w3987 = (~pi0633 & ~w2402) | (~pi0633 & w10178) | (~w2402 & w10178);
assign w3988 = ~w3986 & ~w3987;
assign w3989 = w3368 & ~w3721;
assign w3990 = (~pi0634 & ~w3367) | (~pi0634 & w10179) | (~w3367 & w10179);
assign w3991 = ~w3989 & ~w3990;
assign w3992 = w2401 & w10180;
assign w3993 = (~pi0635 & ~w2401) | (~pi0635 & w10181) | (~w2401 & w10181);
assign w3994 = pi1150 & ~w3992;
assign w3995 = ~w3993 & w3994;
assign w3996 = w2400 & w10182;
assign w3997 = pi0636 & ~w3996;
assign w3998 = w3368 & ~w3713;
assign w3999 = (~pi0637 & ~w3367) | (~pi0637 & w10183) | (~w3367 & w10183);
assign w4000 = ~w3998 & ~w3999;
assign w4001 = w2445 & ~w2624;
assign w4002 = (~pi0638 & ~w2402) | (~pi0638 & w10184) | (~w2402 & w10184);
assign w4003 = ~w4001 & ~w4002;
assign w4004 = pi0192 & w3435;
assign w4005 = pi0207 & w3369;
assign w4006 = pi1924 & w3363;
assign w4007 = ~w4004 & ~w4005;
assign w4008 = ~w4006 & w4007;
assign w4009 = w3376 & ~w4008;
assign w4010 = (~pi0639 & ~w3367) | (~pi0639 & w10185) | (~w3367 & w10185);
assign w4011 = ~w4009 & ~w4010;
assign w4012 = pi0479 & w3435;
assign w4013 = pi0866 & w3369;
assign w4014 = pi0820 & w3363;
assign w4015 = ~w4012 & ~w4013;
assign w4016 = ~w4014 & w4015;
assign w4017 = w3368 & ~w4016;
assign w4018 = (~pi0641 & ~w3367) | (~pi0641 & w10186) | (~w3367 & w10186);
assign w4019 = ~w4017 & ~w4018;
assign w4020 = pi0857 & w3383;
assign w4021 = pi1933 & w3481;
assign w4022 = pi1157 & ~pi1158;
assign w4023 = pi1883 & w4022;
assign w4024 = ~w4020 & ~w4021;
assign w4025 = ~w4023 & w4024;
assign w4026 = w3480 & ~w4025;
assign w4027 = (~pi0642 & ~w3387) | (~pi0642 & w10187) | (~w3387 & w10187);
assign w4028 = ~w4026 & ~w4027;
assign w4029 = w3387 & w10189;
assign w4030 = (w3387 & w10190) | (w3387 & w10191) | (w10190 & w10191);
assign w4031 = ~w4029 & w4030;
assign w4032 = pi0883 & w4022;
assign w4033 = pi0951 & w3481;
assign w4034 = pi0858 & w3383;
assign w4035 = ~w4032 & ~w4033;
assign w4036 = ~w4034 & w4035;
assign w4037 = w3480 & ~w4036;
assign w4038 = (~pi0644 & ~w3387) | (~pi0644 & w10192) | (~w3387 & w10192);
assign w4039 = ~w4037 & ~w4038;
assign w4040 = pi0828 & w3363;
assign w4041 = pi0882 & w3435;
assign w4042 = pi0950 & w3369;
assign w4043 = ~w4040 & ~w4041;
assign w4044 = ~w4042 & w4043;
assign w4045 = w3434 & ~w4044;
assign w4046 = (~pi0645 & ~w3367) | (~pi0645 & w10193) | (~w3367 & w10193);
assign w4047 = ~w4045 & ~w4046;
assign w4048 = pi1933 & w4022;
assign w4049 = pi1958 & w3481;
assign w4050 = pi0854 & w3383;
assign w4051 = ~w4048 & ~w4049;
assign w4052 = ~w4050 & w4051;
assign w4053 = w3480 & ~w4052;
assign w4054 = (~pi0646 & ~w3387) | (~pi0646 & w10194) | (~w3387 & w10194);
assign w4055 = ~w4053 & ~w4054;
assign w4056 = w3387 & w10196;
assign w4057 = (~pi0647 & ~w3387) | (~pi0647 & w10197) | (~w3387 & w10197);
assign w4058 = ~w4056 & ~w4057;
assign w4059 = w3434 & ~w3729;
assign w4060 = (~pi0648 & ~w3367) | (~pi0648 & w10198) | (~w3367 & w10198);
assign w4061 = ~w4059 & ~w4060;
assign w4062 = pi0191 & w4022;
assign w4063 = pi0206 & w3481;
assign w4064 = pi1925 & w3383;
assign w4065 = ~w4062 & ~w4063;
assign w4066 = ~w4064 & w4065;
assign w4067 = w3480 & ~w4066;
assign w4068 = (~pi0649 & ~w3387) | (~pi0649 & w10199) | (~w3387 & w10199);
assign w4069 = ~w4067 & ~w4068;
assign w4070 = pi0231 & w4022;
assign w4071 = pi0481 & w3481;
assign w4072 = pi0851 & w3383;
assign w4073 = ~w4070 & ~w4071;
assign w4074 = ~w4072 & w4073;
assign w4075 = w3480 & ~w4074;
assign w4076 = (~pi0650 & ~w3387) | (~pi0650 & w10200) | (~w3387 & w10200);
assign w4077 = ~w4075 & ~w4076;
assign w4078 = w3434 & ~w3713;
assign w4079 = (~pi0651 & ~w3367) | (~pi0651 & w10201) | (~w3367 & w10201);
assign w4080 = ~w4078 & ~w4079;
assign w4081 = pi0207 & w3435;
assign w4082 = pi0235 & w3369;
assign w4083 = pi0833 & w3363;
assign w4084 = ~w4081 & ~w4082;
assign w4085 = ~w4083 & w4084;
assign w4086 = w3434 & ~w4085;
assign w4087 = (~pi0652 & ~w3367) | (~pi0652 & w10202) | (~w3367 & w10202);
assign w4088 = ~w4086 & ~w4087;
assign w4089 = w3434 & ~w3896;
assign w4090 = (~pi0653 & ~w3367) | (~pi0653 & w10203) | (~w3367 & w10203);
assign w4091 = ~w4089 & ~w4090;
assign w4092 = pi0832 & w3363;
assign w4093 = pi0882 & w3369;
assign w4094 = pi0819 & w3435;
assign w4095 = ~w4092 & ~w4093;
assign w4096 = ~w4094 & w4095;
assign w4097 = w3434 & ~w4096;
assign w4098 = (~pi0654 & ~w3367) | (~pi0654 & w10204) | (~w3367 & w10204);
assign w4099 = ~w4097 & ~w4098;
assign w4100 = w3376 & ~w4044;
assign w4101 = (~pi0655 & ~w3367) | (~pi0655 & w10205) | (~w3367 & w10205);
assign w4102 = ~w4100 & ~w4101;
assign w4103 = w3367 & w10206;
assign w4104 = (~pi0656 & ~w3367) | (~pi0656 & w10207) | (~w3367 & w10207);
assign w4105 = ~w4103 & ~w4104;
assign w4106 = w2400 & w10208;
assign w4107 = pi0657 & ~w4106;
assign w4108 = pi0814 & w4106;
assign w4109 = ~w4107 & ~w4108;
assign w4110 = pi0333 & w4022;
assign w4111 = pi0818 & w3481;
assign w4112 = pi0850 & w3383;
assign w4113 = ~w4110 & ~w4111;
assign w4114 = ~w4112 & w4113;
assign w4115 = w3401 & ~w4114;
assign w4116 = (~pi0658 & ~w3387) | (~pi0658 & w10209) | (~w3387 & w10209);
assign w4117 = ~w4115 & ~w4116;
assign w4118 = w3376 & ~w3896;
assign w4119 = (~pi0659 & ~w3367) | (~pi0659 & w10210) | (~w3367 & w10210);
assign w4120 = ~w4118 & ~w4119;
assign w4121 = w3376 & ~w3440;
assign w4122 = (~pi0660 & ~w3367) | (~pi0660 & w10211) | (~w3367 & w10211);
assign w4123 = ~w4121 & ~w4122;
assign w4124 = w3388 & ~w4025;
assign w4125 = (~pi0661 & ~w3387) | (~pi0661 & w10212) | (~w3387 & w10212);
assign w4126 = ~w4124 & ~w4125;
assign w4127 = pi1981 & w4022;
assign w4128 = pi1959 & w3481;
assign w4129 = pi0853 & w3383;
assign w4130 = ~w4127 & ~w4128;
assign w4131 = ~w4129 & w4130;
assign w4132 = w3388 & ~w4131;
assign w4133 = (~pi0662 & ~w3387) | (~pi0662 & w10213) | (~w3387 & w10213);
assign w4134 = ~w4132 & ~w4133;
assign w4135 = pi0206 & w4022;
assign w4136 = pi0231 & w3481;
assign w4137 = pi0852 & w3383;
assign w4138 = ~w4135 & ~w4136;
assign w4139 = ~w4137 & w4138;
assign w4140 = w3388 & ~w4139;
assign w4141 = (~pi0663 & ~w3387) | (~pi0663 & w10214) | (~w3387 & w10214);
assign w4142 = ~w4140 & ~w4141;
assign w4143 = pi1853 & w4022;
assign w4144 = pi1925 & w3481;
assign w4145 = pi0855 & w3383;
assign w4146 = ~w4143 & ~w4144;
assign w4147 = ~w4145 & w4146;
assign w4148 = w3401 & ~w4147;
assign w4149 = (~pi0664 & ~w3387) | (~pi0664 & w10215) | (~w3387 & w10215);
assign w4150 = ~w4148 & ~w4149;
assign w4151 = w3401 & ~w4052;
assign w4152 = (~pi0665 & ~w3387) | (~pi0665 & w10216) | (~w3387 & w10216);
assign w4153 = ~w4151 & ~w4152;
assign w4154 = w3434 & ~w3745;
assign w4155 = (~pi0666 & ~w3367) | (~pi0666 & w10217) | (~w3367 & w10217);
assign w4156 = ~w4154 & ~w4155;
assign w4157 = w3421 & ~w3440;
assign w4158 = (~pi0667 & ~w3367) | (~pi0667 & w10218) | (~w3367 & w10218);
assign w4159 = ~w4157 & ~w4158;
assign w4160 = w3421 & ~w4016;
assign w4161 = (~pi0668 & ~w3367) | (~pi0668 & w10219) | (~w3367 & w10219);
assign w4162 = ~w4160 & ~w4161;
assign w4163 = w3421 & ~w3904;
assign w4164 = (~pi0669 & ~w3367) | (~pi0669 & w10220) | (~w3367 & w10220);
assign w4165 = ~w4163 & ~w4164;
assign w4166 = w3421 & ~w3896;
assign w4167 = (~pi0670 & ~w3367) | (~pi0670 & w10221) | (~w3367 & w10221);
assign w4168 = ~w4166 & ~w4167;
assign w4169 = pi0212 & w3435;
assign w4170 = pi0334 & w3369;
assign w4171 = pi0834 & w3363;
assign w4172 = ~w4169 & ~w4170;
assign w4173 = ~w4171 & w4172;
assign w4174 = w3421 & ~w4173;
assign w4175 = (~pi0671 & ~w3367) | (~pi0671 & w10222) | (~w3367 & w10222);
assign w4176 = ~w4174 & ~w4175;
assign w4177 = w3421 & ~w4085;
assign w4178 = (~pi0672 & ~w3367) | (~pi0672 & w10223) | (~w3367 & w10223);
assign w4179 = ~w4177 & ~w4178;
assign w4180 = pi0196 & w3435;
assign w4181 = pi0212 & w3369;
assign w4182 = pi1934 & w3363;
assign w4183 = ~w4180 & ~w4181;
assign w4184 = ~w4182 & w4183;
assign w4185 = w3421 & ~w4184;
assign w4186 = (~pi0673 & ~w3367) | (~pi0673 & w10224) | (~w3367 & w10224);
assign w4187 = ~w4185 & ~w4186;
assign w4188 = w3421 & ~w4096;
assign w4189 = (~pi0674 & ~w3367) | (~pi0674 & w10225) | (~w3367 & w10225);
assign w4190 = ~w4188 & ~w4189;
assign w4191 = pi1958 & w4022;
assign w4192 = pi1947 & w3481;
assign w4193 = pi0848 & w3383;
assign w4194 = ~w4191 & ~w4192;
assign w4195 = ~w4193 & w4194;
assign w4196 = w3411 & ~w4195;
assign w4197 = (~pi0675 & ~w3387) | (~pi0675 & w10226) | (~w3387 & w10226);
assign w4198 = ~w4196 & ~w4197;
assign w4199 = pi0846 & w3383;
assign w4200 = pi0883 & w3481;
assign w4201 = pi0818 & w4022;
assign w4202 = ~w4199 & ~w4200;
assign w4203 = ~w4201 & w4202;
assign w4204 = w3411 & ~w4203;
assign w4205 = (~pi0676 & ~w3387) | (~pi0676 & w10227) | (~w3387 & w10227);
assign w4206 = ~w4204 & ~w4205;
assign w4207 = w3411 & ~w4114;
assign w4208 = (~pi0677 & ~w3387) | (~pi0677 & w10228) | (~w3387 & w10228);
assign w4209 = ~w4207 & ~w4208;
assign w4210 = w3411 & ~w4074;
assign w4211 = (~pi0678 & ~w3387) | (~pi0678 & w10229) | (~w3387 & w10229);
assign w4212 = ~w4210 & ~w4211;
assign w4213 = pi0847 & w3383;
assign w4214 = pi0211 & w4022;
assign w4215 = pi0333 & w3481;
assign w4216 = ~w4213 & ~w4214;
assign w4217 = ~w4215 & w4216;
assign w4218 = w3411 & ~w4217;
assign w4219 = (~pi0679 & ~w3387) | (~pi0679 & w10230) | (~w3387 & w10230);
assign w4220 = ~w4218 & ~w4219;
assign w4221 = pi1933 & w3383;
assign w4222 = pi0211 & w3481;
assign w4223 = pi0195 & w4022;
assign w4224 = ~w4221 & ~w4222;
assign w4225 = ~w4223 & w4224;
assign w4226 = w3411 & ~w4225;
assign w4227 = (~pi0680 & ~w3387) | (~pi0680 & w10231) | (~w3387 & w10231);
assign w4228 = ~w4226 & ~w4227;
assign w4229 = w3411 & ~w4066;
assign w4230 = (~pi0681 & ~w3387) | (~pi0681 & w10232) | (~w3387 & w10232);
assign w4231 = ~w4229 & ~w4230;
assign w4232 = w3411 & ~w4131;
assign w4233 = (~pi0682 & ~w3387) | (~pi0682 & w10233) | (~w3387 & w10233);
assign w4234 = ~w4232 & ~w4233;
assign w4235 = w3411 & ~w4052;
assign w4236 = (~pi0683 & ~w3387) | (~pi0683 & w10234) | (~w3387 & w10234);
assign w4237 = ~w4235 & ~w4236;
assign w4238 = pi1925 & w4022;
assign w4239 = pi1981 & w3481;
assign w4240 = pi0845 & w3383;
assign w4241 = ~w4238 & ~w4239;
assign w4242 = ~w4240 & w4241;
assign w4243 = w3411 & ~w4242;
assign w4244 = (~pi0684 & ~w3387) | (~pi0684 & w10235) | (~w3387 & w10235);
assign w4245 = ~w4243 & ~w4244;
assign w4246 = w3411 & ~w4025;
assign w4247 = (~pi0685 & ~w3387) | (~pi0685 & w10236) | (~w3387 & w10236);
assign w4248 = ~w4246 & ~w4247;
assign w4249 = w3411 & ~w4147;
assign w4250 = (~pi0686 & ~w3387) | (~pi0686 & w10237) | (~w3387 & w10237);
assign w4251 = ~w4249 & ~w4250;
assign w4252 = pi0951 & w4022;
assign w4253 = pi1883 & w3481;
assign w4254 = pi0856 & w3383;
assign w4255 = ~w4252 & ~w4253;
assign w4256 = ~w4254 & w4255;
assign w4257 = w3411 & ~w4256;
assign w4258 = (~pi0687 & ~w3387) | (~pi0687 & w10238) | (~w3387 & w10238);
assign w4259 = ~w4257 & ~w4258;
assign w4260 = pi0916 & w4022;
assign w4261 = pi1853 & w3481;
assign w4262 = pi0859 & w3383;
assign w4263 = ~w4260 & ~w4261;
assign w4264 = ~w4262 & w4263;
assign w4265 = w3411 & ~w4264;
assign w4266 = (~pi0688 & ~w3387) | (~pi0688 & w10239) | (~w3387 & w10239);
assign w4267 = ~w4265 & ~w4266;
assign w4268 = w3411 & ~w4036;
assign w4269 = (~pi0689 & ~w3387) | (~pi0689 & w10240) | (~w3387 & w10240);
assign w4270 = ~w4268 & ~w4269;
assign w4271 = w3401 & ~w4195;
assign w4272 = (~pi0690 & ~w3387) | (~pi0690 & w10241) | (~w3387 & w10241);
assign w4273 = ~w4271 & ~w4272;
assign w4274 = w3401 & ~w4203;
assign w4275 = (~pi0691 & ~w3387) | (~pi0691 & w10242) | (~w3387 & w10242);
assign w4276 = ~w4274 & ~w4275;
assign w4277 = pi0481 & w4022;
assign w4278 = pi0870 & w3481;
assign w4279 = pi0849 & w3383;
assign w4280 = ~w4277 & ~w4278;
assign w4281 = ~w4279 & w4280;
assign w4282 = w3401 & ~w4281;
assign w4283 = (~pi0692 & ~w3387) | (~pi0692 & w10243) | (~w3387 & w10243);
assign w4284 = ~w4282 & ~w4283;
assign w4285 = w3401 & ~w4217;
assign w4286 = (~pi0693 & ~w3387) | (~pi0693 & w10244) | (~w3387 & w10244);
assign w4287 = ~w4285 & ~w4286;
assign w4288 = w3401 & ~w4139;
assign w4289 = (~pi0694 & ~w3387) | (~pi0694 & w10245) | (~w3387 & w10245);
assign w4290 = ~w4288 & ~w4289;
assign w4291 = w3401 & ~w4225;
assign w4292 = (~pi0695 & ~w3387) | (~pi0695 & w10246) | (~w3387 & w10246);
assign w4293 = ~w4291 & ~w4292;
assign w4294 = w3401 & ~w4066;
assign w4295 = (~pi0696 & ~w3387) | (~pi0696 & w10247) | (~w3387 & w10247);
assign w4296 = ~w4294 & ~w4295;
assign w4297 = w3401 & ~w4131;
assign w4298 = (~pi0697 & ~w3387) | (~pi0697 & w10248) | (~w3387 & w10248);
assign w4299 = ~w4297 & ~w4298;
assign w4300 = w3421 & ~w3737;
assign w4301 = (~pi0698 & ~w3367) | (~pi0698 & w10249) | (~w3367 & w10249);
assign w4302 = ~w4300 & ~w4301;
assign w4303 = w3401 & ~w4242;
assign w4304 = (~pi0699 & ~w3387) | (~pi0699 & w10250) | (~w3387 & w10250);
assign w4305 = ~w4303 & ~w4304;
assign w4306 = pi1886 & w3435;
assign w4307 = pi1934 & w3369;
assign w4308 = pi0826 & w3363;
assign w4309 = ~w4306 & ~w4307;
assign w4310 = ~w4308 & w4309;
assign w4311 = w3421 & ~w4310;
assign w4312 = (~pi0700 & ~w3367) | (~pi0700 & w10251) | (~w3367 & w10251);
assign w4313 = ~w4311 & ~w4312;
assign w4314 = w3401 & ~w4025;
assign w4315 = (~pi0701 & ~w3387) | (~pi0701 & w10252) | (~w3387 & w10252);
assign w4316 = ~w4314 & ~w4315;
assign w4317 = w3401 & ~w4256;
assign w4318 = (~pi0702 & ~w3387) | (~pi0702 & w10253) | (~w3387 & w10253);
assign w4319 = ~w4317 & ~w4318;
assign w4320 = w3401 & ~w4264;
assign w4321 = (~pi0703 & ~w3387) | (~pi0703 & w10254) | (~w3387 & w10254);
assign w4322 = ~w4320 & ~w4321;
assign w4323 = w3401 & ~w4036;
assign w4324 = (~pi0704 & ~w3387) | (~pi0704 & w10255) | (~w3387 & w10255);
assign w4325 = ~w4323 & ~w4324;
assign w4326 = w3388 & ~w4195;
assign w4327 = (~pi0705 & ~w3387) | (~pi0705 & w10256) | (~w3387 & w10256);
assign w4328 = ~w4326 & ~w4327;
assign w4329 = w3388 & ~w4203;
assign w4330 = (~pi0706 & ~w3387) | (~pi0706 & w10257) | (~w3387 & w10257);
assign w4331 = ~w4329 & ~w4330;
assign w4332 = w3388 & ~w4281;
assign w4333 = (~pi0707 & ~w3387) | (~pi0707 & w10258) | (~w3387 & w10258);
assign w4334 = ~w4332 & ~w4333;
assign w4335 = w3388 & ~w4114;
assign w4336 = (~pi0708 & ~w3387) | (~pi0708 & w10259) | (~w3387 & w10259);
assign w4337 = ~w4335 & ~w4336;
assign w4338 = w3388 & ~w4074;
assign w4339 = (~pi0709 & ~w3387) | (~pi0709 & w10260) | (~w3387 & w10260);
assign w4340 = ~w4338 & ~w4339;
assign w4341 = w3388 & ~w4217;
assign w4342 = (~pi0710 & ~w3387) | (~pi0710 & w10261) | (~w3387 & w10261);
assign w4343 = ~w4341 & ~w4342;
assign w4344 = w3401 & ~w4074;
assign w4345 = (~pi0711 & ~w3387) | (~pi0711 & w10262) | (~w3387 & w10262);
assign w4346 = ~w4344 & ~w4345;
assign w4347 = w3388 & ~w4225;
assign w4348 = (~pi0712 & ~w3387) | (~pi0712 & w10263) | (~w3387 & w10263);
assign w4349 = ~w4347 & ~w4348;
assign w4350 = w3388 & ~w4066;
assign w4351 = (~pi0713 & ~w3387) | (~pi0713 & w10264) | (~w3387 & w10264);
assign w4352 = ~w4350 & ~w4351;
assign w4353 = pi0915 & w3435;
assign w4354 = pi1852 & w3369;
assign w4355 = pi0830 & w3363;
assign w4356 = ~w4353 & ~w4354;
assign w4357 = ~w4355 & w4356;
assign w4358 = w3421 & ~w4357;
assign w4359 = (~pi0714 & ~w3367) | (~pi0714 & w10265) | (~w3367 & w10265);
assign w4360 = ~w4358 & ~w4359;
assign w4361 = w3388 & ~w4052;
assign w4362 = (~pi0715 & ~w3387) | (~pi0715 & w10266) | (~w3387 & w10266);
assign w4363 = ~w4361 & ~w4362;
assign w4364 = w3388 & ~w4242;
assign w4365 = (~pi0716 & ~w3387) | (~pi0716 & w10267) | (~w3387 & w10267);
assign w4366 = ~w4364 & ~w4365;
assign w4367 = w3388 & ~w4147;
assign w4368 = (~pi0717 & ~w3387) | (~pi0717 & w10268) | (~w3387 & w10268);
assign w4369 = ~w4367 & ~w4368;
assign w4370 = w3388 & ~w4256;
assign w4371 = (~pi0718 & ~w3387) | (~pi0718 & w10269) | (~w3387 & w10269);
assign w4372 = ~w4370 & ~w4371;
assign w4373 = w3388 & ~w4264;
assign w4374 = (~pi0719 & ~w3387) | (~pi0719 & w10270) | (~w3387 & w10270);
assign w4375 = ~w4373 & ~w4374;
assign w4376 = w3421 & ~w4044;
assign w4377 = (~pi0720 & ~w3367) | (~pi0720 & w10271) | (~w3367 & w10271);
assign w4378 = ~w4376 & ~w4377;
assign w4379 = pi0870 & w4022;
assign w4380 = pi0916 & w3481;
assign w4381 = pi0844 & w3383;
assign w4382 = ~w4379 & ~w4380;
assign w4383 = ~w4381 & w4382;
assign w4384 = w3388 & ~w4383;
assign w4385 = (~pi0721 & ~w3387) | (~pi0721 & w10272) | (~w3387 & w10272);
assign w4386 = ~w4384 & ~w4385;
assign w4387 = w3388 & ~w4036;
assign w4388 = (~pi0722 & ~w3387) | (~pi0722 & w10273) | (~w3387 & w10273);
assign w4389 = ~w4387 & ~w4388;
assign w4390 = w3376 & ~w4096;
assign w4391 = (~pi0723 & ~w3367) | (~pi0723 & w10274) | (~w3367 & w10274);
assign w4392 = ~w4390 & ~w4391;
assign w4393 = w3376 & ~w4016;
assign w4394 = (~pi0724 & ~w3367) | (~pi0724 & w10275) | (~w3367 & w10275);
assign w4395 = ~w4393 & ~w4394;
assign w4396 = w3376 & ~w3904;
assign w4397 = (~pi0725 & ~w3367) | (~pi0725 & w10276) | (~w3367 & w10276);
assign w4398 = ~w4396 & ~w4397;
assign w4399 = w3376 & ~w4173;
assign w4400 = (~pi0726 & ~w3367) | (~pi0726 & w10277) | (~w3367 & w10277);
assign w4401 = ~w4399 & ~w4400;
assign w4402 = w3376 & ~w4085;
assign w4403 = (~pi0727 & ~w3367) | (~pi0727 & w10278) | (~w3367 & w10278);
assign w4404 = ~w4402 & ~w4403;
assign w4405 = w3376 & ~w4184;
assign w4406 = (~pi0728 & ~w3367) | (~pi0728 & w10279) | (~w3367 & w10279);
assign w4407 = ~w4405 & ~w4406;
assign w4408 = w3376 & ~w3713;
assign w4409 = (~pi0729 & ~w3367) | (~pi0729 & w10280) | (~w3367 & w10280);
assign w4410 = ~w4408 & ~w4409;
assign w4411 = w3376 & ~w4310;
assign w4412 = (~pi0730 & ~w3367) | (~pi0730 & w10281) | (~w3367 & w10281);
assign w4413 = ~w4411 & ~w4412;
assign w4414 = w3376 & ~w3721;
assign w4415 = (~pi0731 & ~w3367) | (~pi0731 & w10282) | (~w3367 & w10282);
assign w4416 = ~w4414 & ~w4415;
assign w4417 = w3376 & ~w3729;
assign w4418 = (~pi0732 & ~w3367) | (~pi0732 & w10283) | (~w3367 & w10283);
assign w4419 = ~w4417 & ~w4418;
assign w4420 = w3376 & ~w4357;
assign w4421 = (~pi0733 & ~w3367) | (~pi0733 & w10284) | (~w3367 & w10284);
assign w4422 = ~w4420 & ~w4421;
assign w4423 = w3434 & ~w4016;
assign w4424 = (~pi0734 & ~w3367) | (~pi0734 & w10285) | (~w3367 & w10285);
assign w4425 = ~w4423 & ~w4424;
assign w4426 = w3434 & ~w3904;
assign w4427 = (~pi0735 & ~w3367) | (~pi0735 & w10286) | (~w3367 & w10286);
assign w4428 = ~w4426 & ~w4427;
assign w4429 = w3434 & ~w4173;
assign w4430 = (~pi0736 & ~w3367) | (~pi0736 & w10287) | (~w3367 & w10287);
assign w4431 = ~w4429 & ~w4430;
assign w4432 = w3434 & ~w4008;
assign w4433 = (~pi0737 & ~w3367) | (~pi0737 & w10288) | (~w3367 & w10288);
assign w4434 = ~w4432 & ~w4433;
assign w4435 = w3434 & ~w4184;
assign w4436 = (~pi0738 & ~w3367) | (~pi0738 & w10289) | (~w3367 & w10289);
assign w4437 = ~w4435 & ~w4436;
assign w4438 = w3411 & ~w4383;
assign w4439 = (~pi0739 & ~w3387) | (~pi0739 & w10290) | (~w3387 & w10290);
assign w4440 = ~w4438 & ~w4439;
assign w4441 = w3434 & ~w3737;
assign w4442 = (~pi0740 & ~w3367) | (~pi0740 & w10291) | (~w3367 & w10291);
assign w4443 = ~w4441 & ~w4442;
assign w4444 = w3434 & ~w4310;
assign w4445 = (~pi0741 & ~w3367) | (~pi0741 & w10292) | (~w3367 & w10292);
assign w4446 = ~w4444 & ~w4445;
assign w4447 = w3434 & ~w3721;
assign w4448 = (~pi0742 & ~w3367) | (~pi0742 & w10293) | (~w3367 & w10293);
assign w4449 = ~w4447 & ~w4448;
assign w4450 = w3434 & ~w3762;
assign w4451 = (~pi0743 & ~w3367) | (~pi0743 & w10294) | (~w3367 & w10294);
assign w4452 = ~w4450 & ~w4451;
assign w4453 = w3421 & ~w3762;
assign w4454 = (~pi0744 & ~w3367) | (~pi0744 & w10295) | (~w3367 & w10295);
assign w4455 = ~w4453 & ~w4454;
assign w4456 = w3434 & ~w4357;
assign w4457 = (~pi0745 & ~w3367) | (~pi0745 & w10296) | (~w3367 & w10296);
assign w4458 = ~w4456 & ~w4457;
assign w4459 = (~pi0746 & ~w3387) | (~pi0746 & w9960) | (~w3387 & w9960);
assign w4460 = (pi1145 & ~w3387) | (pi1145 & w10297) | (~w3387 & w10297);
assign w4461 = ~w4459 & w4460;
assign w4462 = w3411 & ~w4139;
assign w4463 = (~pi0747 & ~w3387) | (~pi0747 & w10298) | (~w3387 & w10298);
assign w4464 = ~w4462 & ~w4463;
assign w4465 = w3411 & ~w4281;
assign w4466 = (~pi0748 & ~w3387) | (~pi0748 & w10299) | (~w3387 & w10299);
assign w4467 = ~w4465 & ~w4466;
assign w4468 = w3421 & ~w4008;
assign w4469 = (~pi0749 & ~w3367) | (~pi0749 & w10300) | (~w3367 & w10300);
assign w4470 = ~w4468 & ~w4469;
assign w4471 = w3367 & w10301;
assign w4472 = (~pi0750 & ~w3367) | (~pi0750 & w10302) | (~w3367 & w10302);
assign w4473 = ~w4471 & ~w4472;
assign w4474 = pi0751 & ~w4106;
assign w4475 = pi0947 & w4106;
assign w4476 = ~w4474 & ~w4475;
assign w4477 = w3368 & ~w4044;
assign w4478 = (~pi0752 & ~w3367) | (~pi0752 & w10303) | (~w3367 & w10303);
assign w4479 = ~w4477 & ~w4478;
assign w4480 = w3368 & ~w4310;
assign w4481 = (~pi0753 & ~w3367) | (~pi0753 & w10304) | (~w3367 & w10304);
assign w4482 = ~w4480 & ~w4481;
assign w4483 = w3480 & ~w4195;
assign w4484 = (~pi0754 & ~w3387) | (~pi0754 & w10305) | (~w3387 & w10305);
assign w4485 = ~w4483 & ~w4484;
assign w4486 = w3480 & ~w4203;
assign w4487 = (~pi0755 & ~w3387) | (~pi0755 & w10306) | (~w3387 & w10306);
assign w4488 = ~w4486 & ~w4487;
assign w4489 = w3480 & ~w4281;
assign w4490 = (~pi0756 & ~w3387) | (~pi0756 & w10307) | (~w3387 & w10307);
assign w4491 = ~w4489 & ~w4490;
assign w4492 = w3480 & ~w4114;
assign w4493 = (~pi0757 & ~w3387) | (~pi0757 & w10308) | (~w3387 & w10308);
assign w4494 = ~w4492 & ~w4493;
assign w4495 = w3480 & ~w4217;
assign w4496 = (~pi0758 & ~w3387) | (~pi0758 & w10309) | (~w3387 & w10309);
assign w4497 = ~w4495 & ~w4496;
assign w4498 = w3480 & ~w4139;
assign w4499 = (~pi0759 & ~w3387) | (~pi0759 & w10310) | (~w3387 & w10310);
assign w4500 = ~w4498 & ~w4499;
assign w4501 = w3480 & ~w4225;
assign w4502 = (~pi0760 & ~w3387) | (~pi0760 & w10311) | (~w3387 & w10311);
assign w4503 = ~w4501 & ~w4502;
assign w4504 = w3480 & ~w4131;
assign w4505 = (~pi0761 & ~w3387) | (~pi0761 & w10312) | (~w3387 & w10312);
assign w4506 = ~w4504 & ~w4505;
assign w4507 = w3387 & w10313;
assign w4508 = (~pi0762 & ~w3387) | (~pi0762 & w10314) | (~w3387 & w10314);
assign w4509 = ~w4507 & ~w4508;
assign w4510 = w3387 & w10315;
assign w4511 = (~pi0763 & ~w3387) | (~pi0763 & w10316) | (~w3387 & w10316);
assign w4512 = ~w4510 & ~w4511;
assign w4513 = w3387 & w10317;
assign w4514 = (~pi0764 & ~w3387) | (~pi0764 & w10318) | (~w3387 & w10318);
assign w4515 = ~w4513 & ~w4514;
assign w4516 = w3387 & w10319;
assign w4517 = (~pi0765 & ~w3387) | (~pi0765 & w10320) | (~w3387 & w10320);
assign w4518 = ~w4516 & ~w4517;
assign w4519 = w3387 & w10321;
assign w4520 = (~pi0766 & ~w3387) | (~pi0766 & w10322) | (~w3387 & w10322);
assign w4521 = ~w4519 & ~w4520;
assign w4522 = w3387 & w10323;
assign w4523 = (~pi0767 & ~w3387) | (~pi0767 & w10324) | (~w3387 & w10324);
assign w4524 = ~w4522 & ~w4523;
assign w4525 = w3387 & w10325;
assign w4526 = (~pi0768 & ~w3387) | (~pi0768 & w10326) | (~w3387 & w10326);
assign w4527 = ~w4525 & ~w4526;
assign w4528 = w3387 & w10327;
assign w4529 = (~pi0769 & ~w3387) | (~pi0769 & w10328) | (~w3387 & w10328);
assign w4530 = ~w4528 & ~w4529;
assign w4531 = w3387 & w10329;
assign w4532 = (~pi0770 & ~w3387) | (~pi0770 & w10330) | (~w3387 & w10330);
assign w4533 = ~w4531 & ~w4532;
assign w4534 = w3387 & w10331;
assign w4535 = (~pi0771 & ~w3387) | (~pi0771 & w10332) | (~w3387 & w10332);
assign w4536 = ~w4534 & ~w4535;
assign w4537 = w3387 & w10333;
assign w4538 = ~pi0772 & ~w3480;
assign w4539 = ~w4537 & ~w4538;
assign w4540 = w3480 & ~w4242;
assign w4541 = (~pi0773 & ~w3387) | (~pi0773 & w10334) | (~w3387 & w10334);
assign w4542 = ~w4540 & ~w4541;
assign w4543 = w3480 & ~w4147;
assign w4544 = (~pi0774 & ~w3387) | (~pi0774 & w10335) | (~w3387 & w10335);
assign w4545 = ~w4543 & ~w4544;
assign w4546 = w3480 & ~w4256;
assign w4547 = (~pi0775 & ~w3387) | (~pi0775 & w10336) | (~w3387 & w10336);
assign w4548 = ~w4546 & ~w4547;
assign w4549 = w3480 & ~w4264;
assign w4550 = (~pi0776 & ~w3387) | (~pi0776 & w10337) | (~w3387 & w10337);
assign w4551 = ~w4549 & ~w4550;
assign w4552 = w3480 & ~w4383;
assign w4553 = (~pi0777 & ~w3387) | (~pi0777 & w10338) | (~w3387 & w10338);
assign w4554 = ~w4552 & ~w4553;
assign w4555 = w3368 & ~w3440;
assign w4556 = (~pi0778 & ~w3367) | (~pi0778 & w10339) | (~w3367 & w10339);
assign w4557 = ~w4555 & ~w4556;
assign w4558 = w3368 & ~w4096;
assign w4559 = (~pi0779 & ~w3367) | (~pi0779 & w10340) | (~w3367 & w10340);
assign w4560 = ~w4558 & ~w4559;
assign w4561 = w3368 & ~w4173;
assign w4562 = (~pi0780 & ~w3367) | (~pi0780 & w10341) | (~w3367 & w10341);
assign w4563 = ~w4561 & ~w4562;
assign w4564 = w3368 & ~w4085;
assign w4565 = (~pi0781 & ~w3367) | (~pi0781 & w10342) | (~w3367 & w10342);
assign w4566 = ~w4564 & ~w4565;
assign w4567 = w3368 & ~w4184;
assign w4568 = (~pi0782 & ~w3367) | (~pi0782 & w10343) | (~w3367 & w10343);
assign w4569 = ~w4567 & ~w4568;
assign w4570 = w3368 & ~w4008;
assign w4571 = (~pi0783 & ~w3367) | (~pi0783 & w10344) | (~w3367 & w10344);
assign w4572 = ~w4570 & ~w4571;
assign w4573 = w3367 & w10345;
assign w4574 = (~pi0784 & ~w3367) | (~pi0784 & w10346) | (~w3367 & w10346);
assign w4575 = ~w4573 & ~w4574;
assign w4576 = w3368 & ~w3737;
assign w4577 = (~pi0785 & ~w3367) | (~pi0785 & w10347) | (~w3367 & w10347);
assign w4578 = ~w4576 & ~w4577;
assign w4579 = w3367 & w10348;
assign w4580 = (~pi0786 & ~w3367) | (~pi0786 & w10349) | (~w3367 & w10349);
assign w4581 = ~w4579 & ~w4580;
assign w4582 = w3368 & ~w3729;
assign w4583 = (~pi0787 & ~w3367) | (~pi0787 & w10350) | (~w3367 & w10350);
assign w4584 = ~w4582 & ~w4583;
assign w4585 = w3368 & ~w4357;
assign w4586 = (~pi0788 & ~w3367) | (~pi0788 & w10351) | (~w3367 & w10351);
assign w4587 = ~w4585 & ~w4586;
assign w4588 = w3368 & ~w3745;
assign w4589 = (~pi0789 & ~w3367) | (~pi0789 & w10352) | (~w3367 & w10352);
assign w4590 = ~w4588 & ~w4589;
assign w4591 = w3366 & w10353;
assign w4592 = (~pi0790 & ~w3366) | (~pi0790 & w10354) | (~w3366 & w10354);
assign w4593 = pi1036 & ~w4591;
assign w4594 = ~w4592 & w4593;
assign w4595 = pi0791 & ~w4106;
assign w4596 = pi1935 & w4106;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = pi0792 & ~w4106;
assign w4599 = pi0335 & w4106;
assign w4600 = ~w4598 & ~w4599;
assign w4601 = pi0793 & ~w4106;
assign w4602 = pi0233 & w4106;
assign w4603 = ~w4601 & ~w4602;
assign w4604 = pi0794 & ~w4106;
assign w4605 = pi0213 & w4106;
assign w4606 = ~w4604 & ~w4605;
assign w4607 = pi0795 & ~w4106;
assign w4608 = pi0208 & w4106;
assign w4609 = ~w4607 & ~w4608;
assign w4610 = pi0796 & ~w4106;
assign w4611 = pi0197 & w4106;
assign w4612 = ~w4610 & ~w4611;
assign w4613 = pi0797 & ~w4106;
assign w4614 = pi0193 & w4106;
assign w4615 = ~w4613 & ~w4614;
assign w4616 = pi0798 & ~w4106;
assign w4617 = pi1926 & w4106;
assign w4618 = ~w4616 & ~w4617;
assign w4619 = pi0799 & ~w4106;
assign w4620 = pi1901 & w4106;
assign w4621 = ~w4619 & ~w4620;
assign w4622 = pi0800 & ~w4106;
assign w4623 = pi1875 & w4106;
assign w4624 = ~w4622 & ~w4623;
assign w4625 = pi0801 & ~w4106;
assign w4626 = pi0923 & w4106;
assign w4627 = ~w4625 & ~w4626;
assign w4628 = pi0802 & ~w4106;
assign w4629 = pi0877 & w4106;
assign w4630 = ~w4628 & ~w4629;
assign w4631 = pi0803 & ~w4106;
assign w4632 = pi0871 & w4106;
assign w4633 = ~w4631 & ~w4632;
assign w4634 = pi0804 & ~w4106;
assign w4635 = pi0480 & w4106;
assign w4636 = ~w4634 & ~w4635;
assign w4637 = w3401 & ~w4383;
assign w4638 = (~pi0805 & ~w3387) | (~pi0805 & w10355) | (~w3387 & w10355);
assign w4639 = ~w4637 & ~w4638;
assign w4640 = w602 & w10356;
assign w4641 = pi0806 & ~w4640;
assign w4642 = w613 & w10357;
assign w4643 = pi0807 & ~w4642;
assign w4644 = w3365 & w10358;
assign w4645 = pi0808 & ~w4644;
assign w4646 = ~pi1144 & pi1905;
assign w4647 = pi0946 & ~pi1930;
assign w4648 = pi0809 & ~w4647;
assign w4649 = ~w4646 & ~w4648;
assign w4650 = (~pi0810 & ~w4647) | (~pi0810 & w10359) | (~w4647 & w10359);
assign w4651 = ~w686 & ~w4650;
assign w4652 = w3367 & w10360;
assign w4653 = ~pi0811 & ~w3368;
assign w4654 = ~w4652 & ~w4653;
assign w4655 = pi0890 & pi2032;
assign w4656 = ~pi0247 & ~pi2032;
assign w4657 = ~w4655 & ~w4656;
assign w4658 = w3365 & w10361;
assign w4659 = pi0813 & ~w4658;
assign w4660 = pi0207 & w4658;
assign w4661 = ~w4659 & ~w4660;
assign w4662 = pi0814 & pi2058;
assign w4663 = pi0891 & ~pi2058;
assign w4664 = ~w4662 & ~w4663;
assign w4665 = ~pi0815 & ~pi0908;
assign w4666 = ~w686 & ~w4665;
assign w4667 = pi0891 & pi2060;
assign w4668 = pi0816 & ~pi2060;
assign w4669 = ~w4667 & ~w4668;
assign w4670 = pi0817 & pi2056;
assign w4671 = pi0891 & ~pi2056;
assign w4672 = ~w4670 & ~w4671;
assign w4673 = pi0818 & pi2059;
assign w4674 = pi0891 & ~pi2059;
assign w4675 = ~w4673 & ~w4674;
assign w4676 = pi0819 & pi2057;
assign w4677 = pi0891 & ~pi2057;
assign w4678 = ~w4676 & ~w4677;
assign w4679 = pi0820 & ~w4658;
assign w4680 = pi0235 & w4658;
assign w4681 = ~w4679 & ~w4680;
assign w4682 = w3386 & w10362;
assign w4683 = (~pi0821 & ~w3386) | (~pi0821 & w10363) | (~w3386 & w10363);
assign w4684 = pi1145 & ~w4682;
assign w4685 = ~w4683 & w4684;
assign w4686 = pi0822 & ~w4658;
assign w4687 = pi0915 & w4658;
assign w4688 = ~w4686 & ~w4687;
assign w4689 = pi0823 & ~w4658;
assign w4690 = pi1852 & w4658;
assign w4691 = ~w4689 & ~w4690;
assign w4692 = pi0824 & ~w4658;
assign w4693 = pi1924 & w4658;
assign w4694 = ~w4692 & ~w4693;
assign w4695 = pi0825 & ~w4658;
assign w4696 = pi1886 & w4658;
assign w4697 = ~w4695 & ~w4696;
assign w4698 = pi0826 & ~w4658;
assign w4699 = pi0950 & w4658;
assign w4700 = ~w4698 & ~w4699;
assign w4701 = pi0827 & ~w4658;
assign w4702 = pi0882 & w4658;
assign w4703 = ~w4701 & ~w4702;
assign w4704 = pi0828 & ~w4658;
assign w4705 = pi0819 & w4658;
assign w4706 = ~w4704 & ~w4705;
assign w4707 = pi0829 & ~w4658;
assign w4708 = pi0479 & w4658;
assign w4709 = ~w4707 & ~w4708;
assign w4710 = pi0830 & ~w4658;
assign w4711 = pi0866 & w4658;
assign w4712 = ~w4710 & ~w4711;
assign w4713 = pi0831 & ~w4658;
assign w4714 = pi1934 & w4658;
assign w4715 = ~w4713 & ~w4714;
assign w4716 = pi0832 & ~w4658;
assign w4717 = pi0334 & w4658;
assign w4718 = ~w4716 & ~w4717;
assign w4719 = pi0833 & ~w4658;
assign w4720 = pi0192 & w4658;
assign w4721 = ~w4719 & ~w4720;
assign w4722 = pi0834 & ~w4658;
assign w4723 = pi0196 & w4658;
assign w4724 = ~w4722 & ~w4723;
assign w4725 = pi0835 & ~w4658;
assign w4726 = pi0212 & w4658;
assign w4727 = ~w4725 & ~w4726;
assign w4728 = ~pi0836 & ~w4647;
assign w4729 = pi0449 & ~w4728;
assign w4730 = pi0449 & w4647;
assign w4731 = pi0860 & pi0873;
assign w4732 = ~pi0837 & ~w4731;
assign w4733 = ~w4730 & ~w4732;
assign w4734 = ~pi0841 & ~pi0928;
assign w4735 = ~w686 & ~w4734;
assign w4736 = ~pi0842 & ~pi0927;
assign w4737 = ~w686 & ~w4736;
assign w4738 = ~pi0843 & ~w3387;
assign w4739 = (pi1145 & ~w3387) | (pi1145 & w10364) | (~w3387 & w10364);
assign w4740 = ~w4738 & w4739;
assign w4741 = w3385 & w10365;
assign w4742 = pi0844 & ~w4741;
assign w4743 = pi0481 & w4741;
assign w4744 = ~w4742 & ~w4743;
assign w4745 = pi0845 & ~w4741;
assign w4746 = pi1853 & w4741;
assign w4747 = ~w4745 & ~w4746;
assign w4748 = pi0846 & ~w4741;
assign w4749 = pi0333 & w4741;
assign w4750 = ~w4748 & ~w4749;
assign w4751 = pi0847 & ~w4741;
assign w4752 = pi0195 & w4741;
assign w4753 = ~w4751 & ~w4752;
assign w4754 = pi0848 & ~w4741;
assign w4755 = pi1933 & w4741;
assign w4756 = ~w4754 & ~w4755;
assign w4757 = pi0849 & ~w4741;
assign w4758 = pi0231 & w4741;
assign w4759 = ~w4757 & ~w4758;
assign w4760 = pi0850 & ~w4741;
assign w4761 = pi0211 & w4741;
assign w4762 = ~w4760 & ~w4761;
assign w4763 = pi0851 & ~w4741;
assign w4764 = pi0206 & w4741;
assign w4765 = ~w4763 & ~w4764;
assign w4766 = pi0852 & ~w4741;
assign w4767 = pi0191 & w4741;
assign w4768 = ~w4766 & ~w4767;
assign w4769 = pi0853 & ~w4741;
assign w4770 = pi1925 & w4741;
assign w4771 = ~w4769 & ~w4770;
assign w4772 = pi0854 & ~w4741;
assign w4773 = pi1883 & w4741;
assign w4774 = ~w4772 & ~w4773;
assign w4775 = pi0855 & ~w4741;
assign w4776 = pi0916 & w4741;
assign w4777 = ~w4775 & ~w4776;
assign w4778 = pi0856 & ~w4741;
assign w4779 = pi0883 & w4741;
assign w4780 = ~w4778 & ~w4779;
assign w4781 = pi0857 & ~w4741;
assign w4782 = pi0951 & w4741;
assign w4783 = ~w4781 & ~w4782;
assign w4784 = pi0858 & ~w4741;
assign w4785 = pi0818 & w4741;
assign w4786 = ~w4784 & ~w4785;
assign w4787 = pi0859 & ~w4741;
assign w4788 = pi0870 & w4741;
assign w4789 = ~w4787 & ~w4788;
assign w4790 = pi0860 & ~pi0873;
assign w4791 = ~pi0837 & w3314;
assign w4792 = ~w4790 & ~w4791;
assign w4793 = ~pi2254 & w2264;
assign w4794 = pi0866 & pi2057;
assign w4795 = pi0925 & ~pi2057;
assign w4796 = ~w4794 & ~w4795;
assign w4797 = pi0925 & pi2060;
assign w4798 = pi0867 & ~pi2060;
assign w4799 = ~w4797 & ~w4798;
assign w4800 = pi0868 & pi2035;
assign w4801 = pi0925 & ~pi2035;
assign w4802 = ~w4800 & ~w4801;
assign w4803 = pi0869 & pi2056;
assign w4804 = pi0925 & ~pi2056;
assign w4805 = ~w4803 & ~w4804;
assign w4806 = pi0870 & pi2059;
assign w4807 = pi0925 & ~pi2059;
assign w4808 = ~w4806 & ~w4807;
assign w4809 = pi0871 & pi2058;
assign w4810 = pi0925 & ~pi2058;
assign w4811 = ~w4809 & ~w4810;
assign w4812 = w3385 & w10366;
assign w4813 = pi0872 & ~w4812;
assign w4814 = pi0860 & w3314;
assign w4815 = ~pi2252 & w2414;
assign w4816 = ~pi2253 & w2424;
assign w4817 = pi0877 & pi2058;
assign w4818 = pi1768 & ~pi2058;
assign w4819 = ~w4817 & ~w4818;
assign w4820 = pi0878 & pi2056;
assign w4821 = pi1768 & ~pi2056;
assign w4822 = ~w4820 & ~w4821;
assign w4823 = ~pi0879 & ~pi1930;
assign w4824 = pi1844 & pi1884;
assign w4825 = pi0232 & ~pi0914;
assign w4826 = pi1839 & w4825;
assign w4827 = ~w4823 & ~w4824;
assign w4828 = w4826 & w4827;
assign w4829 = ~w645 & ~w4828;
assign w4830 = pi1879 & pi2134;
assign w4831 = ~pi0880 & ~w4830;
assign w4832 = ~pi1956 & pi1990;
assign w4833 = pi2001 & ~pi2003;
assign w4834 = w4832 & w4833;
assign w4835 = ~w4831 & ~w4834;
assign w4836 = pi0881 & pi2035;
assign w4837 = pi1768 & ~pi2035;
assign w4838 = ~w4836 & ~w4837;
assign w4839 = pi0882 & pi2057;
assign w4840 = pi1768 & ~pi2057;
assign w4841 = ~w4839 & ~w4840;
assign w4842 = pi0883 & pi2059;
assign w4843 = pi1768 & ~pi2059;
assign w4844 = ~w4842 & ~w4843;
assign w4845 = ~pi0884 & ~pi1930;
assign w4846 = pi0868 & pi1172;
assign w4847 = pi0232 & ~pi0909;
assign w4848 = pi1164 & w4847;
assign w4849 = ~w4845 & ~w4846;
assign w4850 = w4848 & w4849;
assign w4851 = ~w629 & ~w4850;
assign w4852 = ~pi0885 & ~pi1930;
assign w4853 = pi0881 & pi1187;
assign w4854 = pi0232 & ~pi0910;
assign w4855 = pi1035 & w4854;
assign w4856 = ~w4852 & ~w4853;
assign w4857 = w4855 & w4856;
assign w4858 = ~w602 & ~w4857;
assign w4859 = ~pi0886 & ~pi1930;
assign w4860 = pi0949 & pi1170;
assign w4861 = pi0232 & ~pi0911;
assign w4862 = pi1169 & w4861;
assign w4863 = ~w4859 & ~w4860;
assign w4864 = w4862 & w4863;
assign w4865 = ~w613 & ~w4864;
assign w4866 = ~pi0887 & ~pi1930;
assign w4867 = pi1177 & pi1850;
assign w4868 = pi0232 & ~pi0907;
assign w4869 = pi1176 & w4868;
assign w4870 = ~w4866 & ~w4867;
assign w4871 = w4869 & w4870;
assign w4872 = ~w637 & ~w4871;
assign w4873 = ~pi0888 & ~pi1930;
assign w4874 = pi1870 & pi1922;
assign w4875 = pi0232 & ~pi0912;
assign w4876 = pi1838 & w4875;
assign w4877 = ~w4873 & ~w4874;
assign w4878 = w4876 & w4877;
assign w4879 = ~w621 & ~w4878;
assign w4880 = ~pi0889 & ~pi1930;
assign w4881 = ~pi0809 & pi1930;
assign w4882 = ~pi0449 & w4881;
assign w4883 = ~w4880 & ~w4882;
assign w4884 = pi1874 & pi2032;
assign w4885 = ~pi0246 & ~pi2032;
assign w4886 = ~w4884 & ~w4885;
assign w4887 = pi0892 & ~pi0893;
assign w4888 = pi0894 & ~pi0895;
assign w4889 = pi0896 & ~pi0897;
assign w4890 = w4888 & w4889;
assign w4891 = w4887 & w4890;
assign w4892 = (pi1878 & ~w4890) | (pi1878 & w10367) | (~w4890 & w10367);
assign w4893 = pi0894 & pi0895;
assign w4894 = pi0893 & w4893;
assign w4895 = w4893 & w10368;
assign w4896 = pi0896 & w4895;
assign w4897 = (~pi0892 & ~w4895) | (~pi0892 & w10369) | (~w4895 & w10369);
assign w4898 = w4895 & w10370;
assign w4899 = w4892 & ~w4897;
assign w4900 = ~w4898 & w4899;
assign w4901 = ~pi0893 & ~w4893;
assign w4902 = ~w4894 & ~w4901;
assign w4903 = w4892 & w4902;
assign w4904 = ~pi0894 & pi1878;
assign w4905 = ~pi0894 & ~pi0895;
assign w4906 = ~w4893 & ~w4905;
assign w4907 = w4892 & w4906;
assign w4908 = ~pi0896 & ~w4895;
assign w4909 = w4892 & ~w4896;
assign w4910 = ~w4908 & w4909;
assign w4911 = (~pi0897 & ~w4893) | (~pi0897 & w10371) | (~w4893 & w10371);
assign w4912 = ~w4895 & ~w4911;
assign w4913 = w4892 & w4912;
assign w4914 = pi2238 & pi2240;
assign w4915 = ~pi2239 & w4914;
assign w4916 = w4914 & w10372;
assign w4917 = pi2241 & ~pi2242;
assign w4918 = w679 & ~w4917;
assign w4919 = w679 & w10373;
assign w4920 = pi2239 & w4914;
assign w4921 = w4917 & w4920;
assign w4922 = w4920 & w10374;
assign w4923 = ~pi2238 & ~pi2239;
assign w4924 = ~pi2240 & w4923;
assign w4925 = ~pi2241 & pi2242;
assign w4926 = ~pi2134 & ~w4925;
assign w4927 = ~pi2104 & w4925;
assign w4928 = w4924 & ~w4926;
assign w4929 = ~w4927 & w4928;
assign w4930 = pi2238 & ~pi2240;
assign w4931 = pi2239 & w4930;
assign w4932 = w4930 & w10375;
assign w4933 = pi2240 & w4923;
assign w4934 = w4923 & w10376;
assign w4935 = ~pi2239 & w4930;
assign w4936 = w4930 & w10377;
assign w4937 = ~pi2240 & w678;
assign w4938 = w678 & w10378;
assign w4939 = w679 & w4917;
assign w4940 = w679 & w10379;
assign w4941 = ~w4916 & ~w4932;
assign w4942 = ~w4934 & ~w4936;
assign w4943 = ~w4938 & w4942;
assign w4944 = ~w4919 & w4941;
assign w4945 = ~w4929 & w10380;
assign w4946 = w4943 & w4944;
assign w4947 = w4945 & w4946;
assign w4948 = pi0221 & ~pi0935;
assign w4949 = ~pi0221 & pi0935;
assign w4950 = ~w4948 & ~w4949;
assign w4951 = pi0225 & ~pi0918;
assign w4952 = ~pi0225 & pi0918;
assign w4953 = pi0217 & ~pi0941;
assign w4954 = ~pi0217 & pi0941;
assign w4955 = ~w4953 & ~w4954;
assign w4956 = ~w4952 & w4955;
assign w4957 = pi1937 & ~w4951;
assign w4958 = ~w4950 & w4957;
assign w4959 = w4956 & w4958;
assign w4960 = pi0899 & ~w4959;
assign w4961 = ~pi0236 & pi0919;
assign w4962 = pi0236 & ~pi0919;
assign w4963 = ~w4961 & ~w4962;
assign w4964 = pi0214 & ~pi0942;
assign w4965 = ~pi0214 & pi0942;
assign w4966 = ~w4964 & ~w4965;
assign w4967 = pi0237 & ~pi0945;
assign w4968 = ~pi0237 & pi0945;
assign w4969 = ~w4967 & ~w4968;
assign w4970 = pi1938 & w4963;
assign w4971 = w4966 & ~w4969;
assign w4972 = w4970 & w4971;
assign w4973 = pi0900 & ~w4972;
assign w4974 = ~pi0226 & pi0922;
assign w4975 = pi0226 & ~pi0922;
assign w4976 = ~w4974 & ~w4975;
assign w4977 = pi0219 & ~pi0944;
assign w4978 = ~pi0219 & pi0944;
assign w4979 = ~w4977 & ~w4978;
assign w4980 = pi0223 & ~pi0937;
assign w4981 = ~pi0223 & pi0937;
assign w4982 = ~w4980 & ~w4981;
assign w4983 = pi1940 & w4976;
assign w4984 = w4979 & ~w4982;
assign w4985 = w4983 & w4984;
assign w4986 = pi0901 & ~w4985;
assign w4987 = ~pi0227 & pi0921;
assign w4988 = pi0227 & ~pi0921;
assign w4989 = ~w4987 & ~w4988;
assign w4990 = pi0218 & ~pi0943;
assign w4991 = ~pi0218 & pi0943;
assign w4992 = ~w4990 & ~w4991;
assign w4993 = pi0222 & ~pi0931;
assign w4994 = ~pi0222 & pi0931;
assign w4995 = ~w4993 & ~w4994;
assign w4996 = pi1936 & w4989;
assign w4997 = w4992 & ~w4995;
assign w4998 = w4996 & w4997;
assign w4999 = pi0902 & ~w4998;
assign w5000 = ~pi0903 & ~pi1930;
assign w5001 = ~w4881 & ~w5000;
assign w5002 = pi0220 & ~pi0934;
assign w5003 = ~pi0220 & pi0934;
assign w5004 = ~w5002 & ~w5003;
assign w5005 = pi0216 & ~pi0940;
assign w5006 = ~pi0216 & pi0940;
assign w5007 = ~w5005 & ~w5006;
assign w5008 = pi0224 & ~pi0917;
assign w5009 = ~pi0224 & pi0917;
assign w5010 = ~w5008 & ~w5009;
assign w5011 = w5007 & w5010;
assign w5012 = pi1941 & ~w5004;
assign w5013 = w5011 & w5012;
assign w5014 = pi0904 & ~w5013;
assign w5015 = pi0239 & ~pi0936;
assign w5016 = ~pi0239 & pi0936;
assign w5017 = ~w5015 & ~w5016;
assign w5018 = pi0238 & ~pi0920;
assign w5019 = ~pi0238 & pi0920;
assign w5020 = pi0215 & ~pi0930;
assign w5021 = ~pi0215 & pi0930;
assign w5022 = ~w5020 & ~w5021;
assign w5023 = ~w5019 & w5022;
assign w5024 = w5022 & w9590;
assign w5025 = pi1939 & ~w5017;
assign w5026 = w5024 & w5025;
assign w5027 = pi0905 & ~w5026;
assign w5028 = pi0906 & pi2056;
assign w5029 = pi1880 & ~pi2056;
assign w5030 = ~w5028 & ~w5029;
assign w5031 = pi0907 & pi1930;
assign w5032 = ~pi1904 & ~pi1930;
assign w5033 = ~w5031 & ~w5032;
assign w5034 = pi0909 & pi1930;
assign w5035 = ~pi1907 & ~pi1930;
assign w5036 = ~w5034 & ~w5035;
assign w5037 = pi0910 & pi1930;
assign w5038 = ~pi1903 & ~pi1930;
assign w5039 = ~w5037 & ~w5038;
assign w5040 = pi0911 & pi1930;
assign w5041 = ~pi1908 & ~pi1930;
assign w5042 = ~w5040 & ~w5041;
assign w5043 = pi0912 & pi1930;
assign w5044 = ~pi1910 & ~pi1930;
assign w5045 = ~w5043 & ~w5044;
assign w5046 = pi1880 & pi2060;
assign w5047 = pi0913 & ~pi2060;
assign w5048 = ~w5046 & ~w5047;
assign w5049 = pi0914 & pi1930;
assign w5050 = ~pi1909 & ~pi1930;
assign w5051 = ~w5049 & ~w5050;
assign w5052 = pi0915 & pi2057;
assign w5053 = pi1880 & ~pi2057;
assign w5054 = ~w5052 & ~w5053;
assign w5055 = pi0916 & pi2059;
assign w5056 = pi1880 & ~pi2059;
assign w5057 = ~w5055 & ~w5056;
assign w5058 = pi0917 & pi1941;
assign w5059 = ~pi0917 & ~pi1941;
assign w5060 = pi1838 & ~w5058;
assign w5061 = ~w5059 & w5060;
assign w5062 = ~pi0918 & pi1937;
assign w5063 = pi0918 & ~pi1937;
assign w5064 = ~w5062 & ~w5063;
assign w5065 = pi1164 & ~w5064;
assign w5066 = pi0919 & pi1938;
assign w5067 = ~pi0919 & ~pi1938;
assign w5068 = pi1035 & ~w5066;
assign w5069 = ~w5067 & w5068;
assign w5070 = ~pi0920 & pi1939;
assign w5071 = pi0920 & ~pi1939;
assign w5072 = ~w5070 & ~w5071;
assign w5073 = pi1169 & ~w5072;
assign w5074 = ~pi0921 & pi1936;
assign w5075 = pi0921 & ~pi1936;
assign w5076 = ~w5074 & ~w5075;
assign w5077 = pi1176 & ~w5076;
assign w5078 = pi0922 & pi1940;
assign w5079 = ~pi0922 & ~pi1940;
assign w5080 = pi1839 & ~w5078;
assign w5081 = ~w5079 & w5080;
assign w5082 = pi0923 & pi2058;
assign w5083 = pi1880 & ~pi2058;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = pi0926 & ~pi0933;
assign w5086 = (~pi0924 & ~w5085) | (~pi0924 & w10381) | (~w5085 & w10381);
assign w5087 = pi1878 & ~w5086;
assign w5088 = w4890 & w10382;
assign w5089 = w5088 & w10384;
assign w5090 = (w5088 & w10385) | (w5088 & w10386) | (w10385 & w10386);
assign w5091 = ~w5089 & w5090;
assign w5092 = ~pi0929 & ~pi1943;
assign w5093 = ~pi0913 & pi1151;
assign w5094 = pi0232 & pi1150;
assign w5095 = ~pi1857 & w5094;
assign w5096 = ~w5092 & ~w5093;
assign w5097 = w5095 & w5096;
assign w5098 = ~w2400 & ~w5097;
assign w5099 = pi0920 & pi1939;
assign w5100 = pi0930 & w5099;
assign w5101 = ~pi0930 & ~w5099;
assign w5102 = (pi1169 & ~w5099) | (pi1169 & w10387) | (~w5099 & w10387);
assign w5103 = ~w5101 & w5102;
assign w5104 = pi0921 & pi1936;
assign w5105 = pi0943 & w5104;
assign w5106 = (~pi0931 & ~w5104) | (~pi0931 & w10388) | (~w5104 & w10388);
assign w5107 = w5104 & w10389;
assign w5108 = pi1176 & ~w5106;
assign w5109 = ~w5107 & w5108;
assign w5110 = w4890 & w10390;
assign w5111 = ~pi0932 & ~w5110;
assign w5112 = pi1878 & ~w5088;
assign w5113 = ~w5111 & w5112;
assign w5114 = ~pi0933 & ~w5088;
assign w5115 = (pi1878 & ~w5088) | (pi1878 & w10391) | (~w5088 & w10391);
assign w5116 = ~w5114 & w5115;
assign w5117 = pi0940 & w5058;
assign w5118 = (~pi0934 & ~w5058) | (~pi0934 & w10392) | (~w5058 & w10392);
assign w5119 = w5058 & w10393;
assign w5120 = pi1838 & ~w5118;
assign w5121 = ~w5119 & w5120;
assign w5122 = pi0918 & pi1937;
assign w5123 = pi0941 & w5122;
assign w5124 = (~pi0935 & ~w5122) | (~pi0935 & w10394) | (~w5122 & w10394);
assign w5125 = w5122 & w10395;
assign w5126 = pi1164 & ~w5124;
assign w5127 = ~w5125 & w5126;
assign w5128 = (~pi0936 & ~w5099) | (~pi0936 & w10396) | (~w5099 & w10396);
assign w5129 = w5099 & w10397;
assign w5130 = pi1169 & ~w5128;
assign w5131 = ~w5129 & w5130;
assign w5132 = pi0944 & w5078;
assign w5133 = (~pi0937 & ~w5078) | (~pi0937 & w10398) | (~w5078 & w10398);
assign w5134 = w5078 & w10399;
assign w5135 = pi1839 & ~w5133;
assign w5136 = ~w5134 & w5135;
assign w5137 = ~pi0938 & pi1931;
assign w5138 = ~pi0816 & pi1153;
assign w5139 = pi0232 & pi1145;
assign w5140 = ~pi1856 & w5139;
assign w5141 = ~w5137 & ~w5138;
assign w5142 = w5140 & w5141;
assign w5143 = ~w3385 & ~w5142;
assign w5144 = ~pi0939 & ~pi1952;
assign w5145 = ~pi0867 & pi1163;
assign w5146 = pi0232 & pi1036;
assign w5147 = ~pi1877 & w5146;
assign w5148 = ~w5144 & ~w5145;
assign w5149 = w5147 & w5148;
assign w5150 = ~w3365 & ~w5149;
assign w5151 = pi0940 & ~w5058;
assign w5152 = ~pi0940 & w5058;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = pi1838 & ~w5153;
assign w5155 = ~pi0941 & ~w5122;
assign w5156 = (pi1164 & ~w5122) | (pi1164 & w10400) | (~w5122 & w10400);
assign w5157 = ~w5155 & w5156;
assign w5158 = pi0942 & ~w5066;
assign w5159 = ~pi0942 & w5066;
assign w5160 = ~w5158 & ~w5159;
assign w5161 = pi1035 & ~w5160;
assign w5162 = ~pi0943 & ~w5104;
assign w5163 = (pi1176 & ~w5104) | (pi1176 & w10401) | (~w5104 & w10401);
assign w5164 = ~w5162 & w5163;
assign w5165 = pi0944 & ~w5078;
assign w5166 = ~pi0944 & w5078;
assign w5167 = ~w5165 & ~w5166;
assign w5168 = pi1839 & ~w5167;
assign w5169 = pi0942 & w5066;
assign w5170 = (~pi0945 & ~w5066) | (~pi0945 & w10402) | (~w5066 & w10402);
assign w5171 = w5066 & w10403;
assign w5172 = pi1035 & ~w5170;
assign w5173 = ~w5171 & w5172;
assign w5174 = pi0947 & pi2058;
assign w5175 = pi1906 & ~pi2058;
assign w5176 = ~w5174 & ~w5175;
assign w5177 = pi0948 & pi2056;
assign w5178 = pi1906 & ~pi2056;
assign w5179 = ~w5177 & ~w5178;
assign w5180 = pi0949 & pi2035;
assign w5181 = pi1906 & ~pi2035;
assign w5182 = ~w5180 & ~w5181;
assign w5183 = pi0950 & pi2057;
assign w5184 = pi1906 & ~pi2057;
assign w5185 = ~w5183 & ~w5184;
assign w5186 = pi0951 & pi2059;
assign w5187 = pi1906 & ~pi2059;
assign w5188 = ~w5186 & ~w5187;
assign w5189 = ~pi0919 & ~pi0942;
assign w5190 = pi1938 & w5189;
assign w5191 = (pi0952 & ~w5189) | (pi0952 & w10404) | (~w5189 & w10404);
assign w5192 = w5189 & w10405;
assign w5193 = ~w5191 & ~w5192;
assign w5194 = (pi0953 & ~w5189) | (pi0953 & w10406) | (~w5189 & w10406);
assign w5195 = w5189 & w10407;
assign w5196 = ~w5194 & ~w5195;
assign w5197 = (pi0954 & ~w5189) | (pi0954 & w10408) | (~w5189 & w10408);
assign w5198 = w5189 & w10409;
assign w5199 = ~w5197 & ~w5198;
assign w5200 = (pi0955 & ~w5189) | (pi0955 & w10410) | (~w5189 & w10410);
assign w5201 = w5189 & w10411;
assign w5202 = ~w5200 & ~w5201;
assign w5203 = (pi0956 & ~w5189) | (pi0956 & w10412) | (~w5189 & w10412);
assign w5204 = w5189 & w10413;
assign w5205 = ~w5203 & ~w5204;
assign w5206 = (pi0957 & ~w5189) | (pi0957 & w10414) | (~w5189 & w10414);
assign w5207 = w5189 & w10415;
assign w5208 = ~w5206 & ~w5207;
assign w5209 = (pi0958 & ~w5189) | (pi0958 & w10416) | (~w5189 & w10416);
assign w5210 = w5189 & w10417;
assign w5211 = ~w5209 & ~w5210;
assign w5212 = (pi0959 & ~w5189) | (pi0959 & w10418) | (~w5189 & w10418);
assign w5213 = w5189 & w10419;
assign w5214 = ~w5212 & ~w5213;
assign w5215 = (pi0960 & ~w5189) | (pi0960 & w10420) | (~w5189 & w10420);
assign w5216 = w5189 & w10421;
assign w5217 = ~w5215 & ~w5216;
assign w5218 = (pi0961 & ~w5189) | (pi0961 & w10422) | (~w5189 & w10422);
assign w5219 = w5189 & w10423;
assign w5220 = ~w5218 & ~w5219;
assign w5221 = ~pi0930 & w5070;
assign w5222 = (pi0962 & ~w5070) | (pi0962 & w10424) | (~w5070 & w10424);
assign w5223 = w5070 & w10425;
assign w5224 = ~w5222 & ~w5223;
assign w5225 = (pi0963 & ~w5070) | (pi0963 & w10426) | (~w5070 & w10426);
assign w5226 = w5070 & w10427;
assign w5227 = ~w5225 & ~w5226;
assign w5228 = (pi0964 & ~w5070) | (pi0964 & w10428) | (~w5070 & w10428);
assign w5229 = w5070 & w10429;
assign w5230 = ~w5228 & ~w5229;
assign w5231 = (pi0965 & ~w5070) | (pi0965 & w10430) | (~w5070 & w10430);
assign w5232 = w5070 & w10431;
assign w5233 = ~w5231 & ~w5232;
assign w5234 = (pi0966 & ~w5070) | (pi0966 & w10432) | (~w5070 & w10432);
assign w5235 = w5070 & w10433;
assign w5236 = ~w5234 & ~w5235;
assign w5237 = (pi0967 & ~w5070) | (pi0967 & w10434) | (~w5070 & w10434);
assign w5238 = w5070 & w10435;
assign w5239 = ~w5237 & ~w5238;
assign w5240 = (pi0968 & ~w5070) | (pi0968 & w10436) | (~w5070 & w10436);
assign w5241 = w5070 & w10437;
assign w5242 = ~w5240 & ~w5241;
assign w5243 = (pi0969 & ~w5070) | (pi0969 & w10438) | (~w5070 & w10438);
assign w5244 = w5070 & w10439;
assign w5245 = ~w5243 & ~w5244;
assign w5246 = (pi0970 & ~w5070) | (pi0970 & w10440) | (~w5070 & w10440);
assign w5247 = w5070 & w10441;
assign w5248 = ~w5246 & ~w5247;
assign w5249 = (pi0971 & ~w5070) | (pi0971 & w10442) | (~w5070 & w10442);
assign w5250 = w5070 & w10443;
assign w5251 = ~w5249 & ~w5250;
assign w5252 = ~pi0943 & w5074;
assign w5253 = (pi0972 & ~w5074) | (pi0972 & w10444) | (~w5074 & w10444);
assign w5254 = w5074 & w10445;
assign w5255 = ~w5253 & ~w5254;
assign w5256 = (pi0973 & ~w5074) | (pi0973 & w10446) | (~w5074 & w10446);
assign w5257 = w5074 & w10447;
assign w5258 = ~w5256 & ~w5257;
assign w5259 = (pi0974 & ~w5074) | (pi0974 & w10448) | (~w5074 & w10448);
assign w5260 = w5074 & w10449;
assign w5261 = ~w5259 & ~w5260;
assign w5262 = (pi0975 & ~w5074) | (pi0975 & w10450) | (~w5074 & w10450);
assign w5263 = w5074 & w10451;
assign w5264 = ~w5262 & ~w5263;
assign w5265 = (pi0976 & ~w5074) | (pi0976 & w10452) | (~w5074 & w10452);
assign w5266 = w5074 & w10453;
assign w5267 = ~w5265 & ~w5266;
assign w5268 = (pi0977 & ~w5074) | (pi0977 & w10454) | (~w5074 & w10454);
assign w5269 = w5074 & w10455;
assign w5270 = ~w5268 & ~w5269;
assign w5271 = (pi0978 & ~w5074) | (pi0978 & w10456) | (~w5074 & w10456);
assign w5272 = w5074 & w10457;
assign w5273 = ~w5271 & ~w5272;
assign w5274 = (pi0979 & ~w5074) | (pi0979 & w10458) | (~w5074 & w10458);
assign w5275 = w5074 & w10459;
assign w5276 = ~w5274 & ~w5275;
assign w5277 = (pi0980 & ~w5074) | (pi0980 & w10460) | (~w5074 & w10460);
assign w5278 = w5074 & w10461;
assign w5279 = ~w5277 & ~w5278;
assign w5280 = (pi0981 & ~w5074) | (pi0981 & w10462) | (~w5074 & w10462);
assign w5281 = w5074 & w10463;
assign w5282 = ~w5280 & ~w5281;
assign w5283 = ~pi0922 & ~pi0944;
assign w5284 = pi1940 & w5283;
assign w5285 = (pi0982 & ~w5283) | (pi0982 & w10464) | (~w5283 & w10464);
assign w5286 = w5283 & w10465;
assign w5287 = ~w5285 & ~w5286;
assign w5288 = (pi0983 & ~w5283) | (pi0983 & w10466) | (~w5283 & w10466);
assign w5289 = w5283 & w10467;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = (pi0984 & ~w5283) | (pi0984 & w10468) | (~w5283 & w10468);
assign w5292 = w5283 & w10469;
assign w5293 = ~w5291 & ~w5292;
assign w5294 = (pi0985 & ~w5283) | (pi0985 & w10470) | (~w5283 & w10470);
assign w5295 = w5283 & w10471;
assign w5296 = ~w5294 & ~w5295;
assign w5297 = (pi0986 & ~w5283) | (pi0986 & w10472) | (~w5283 & w10472);
assign w5298 = w5283 & w10473;
assign w5299 = ~w5297 & ~w5298;
assign w5300 = (pi0987 & ~w5283) | (pi0987 & w10474) | (~w5283 & w10474);
assign w5301 = w5283 & w10475;
assign w5302 = ~w5300 & ~w5301;
assign w5303 = (pi0988 & ~w5283) | (pi0988 & w10476) | (~w5283 & w10476);
assign w5304 = w5283 & w10477;
assign w5305 = ~w5303 & ~w5304;
assign w5306 = (pi0989 & ~w5283) | (pi0989 & w10478) | (~w5283 & w10478);
assign w5307 = w5283 & w10479;
assign w5308 = ~w5306 & ~w5307;
assign w5309 = (pi0990 & ~w5283) | (pi0990 & w10480) | (~w5283 & w10480);
assign w5310 = w5283 & w10481;
assign w5311 = ~w5309 & ~w5310;
assign w5312 = (pi0991 & ~w5283) | (pi0991 & w10482) | (~w5283 & w10482);
assign w5313 = w5283 & w10483;
assign w5314 = ~w5312 & ~w5313;
assign w5315 = ~pi0941 & w5062;
assign w5316 = (pi0992 & ~w5062) | (pi0992 & w10484) | (~w5062 & w10484);
assign w5317 = w5062 & w10485;
assign w5318 = ~w5316 & ~w5317;
assign w5319 = (pi0993 & ~w5062) | (pi0993 & w10486) | (~w5062 & w10486);
assign w5320 = w5062 & w10487;
assign w5321 = ~w5319 & ~w5320;
assign w5322 = (pi0994 & ~w5062) | (pi0994 & w10488) | (~w5062 & w10488);
assign w5323 = w5062 & w10489;
assign w5324 = ~w5322 & ~w5323;
assign w5325 = ~pi0917 & ~pi0940;
assign w5326 = pi1941 & w5325;
assign w5327 = (pi0995 & ~w5325) | (pi0995 & w10490) | (~w5325 & w10490);
assign w5328 = w5325 & w10491;
assign w5329 = ~w5327 & ~w5328;
assign w5330 = (pi0996 & ~w5325) | (pi0996 & w10492) | (~w5325 & w10492);
assign w5331 = w5325 & w10493;
assign w5332 = ~w5330 & ~w5331;
assign w5333 = (pi0997 & ~w5325) | (pi0997 & w10494) | (~w5325 & w10494);
assign w5334 = w5325 & w10495;
assign w5335 = ~w5333 & ~w5334;
assign w5336 = (pi0998 & ~w5325) | (pi0998 & w10496) | (~w5325 & w10496);
assign w5337 = w5325 & w10497;
assign w5338 = ~w5336 & ~w5337;
assign w5339 = (pi0999 & ~w5062) | (pi0999 & w10498) | (~w5062 & w10498);
assign w5340 = w5062 & w10499;
assign w5341 = ~w5339 & ~w5340;
assign w5342 = (pi1000 & ~w5062) | (pi1000 & w10500) | (~w5062 & w10500);
assign w5343 = w5062 & w10501;
assign w5344 = ~w5342 & ~w5343;
assign w5345 = (pi1001 & ~w5325) | (pi1001 & w10502) | (~w5325 & w10502);
assign w5346 = w5325 & w10503;
assign w5347 = ~w5345 & ~w5346;
assign w5348 = (pi1002 & ~w5325) | (pi1002 & w10504) | (~w5325 & w10504);
assign w5349 = w5325 & w10505;
assign w5350 = ~w5348 & ~w5349;
assign w5351 = (pi1003 & ~w5325) | (pi1003 & w10506) | (~w5325 & w10506);
assign w5352 = w5325 & w10507;
assign w5353 = ~w5351 & ~w5352;
assign w5354 = (pi1004 & ~w5325) | (pi1004 & w10508) | (~w5325 & w10508);
assign w5355 = w5325 & w10509;
assign w5356 = ~w5354 & ~w5355;
assign w5357 = (pi1005 & ~w5062) | (pi1005 & w10510) | (~w5062 & w10510);
assign w5358 = w5062 & w10511;
assign w5359 = ~w5357 & ~w5358;
assign w5360 = (pi1006 & ~w5325) | (pi1006 & w10512) | (~w5325 & w10512);
assign w5361 = w5325 & w10513;
assign w5362 = ~w5360 & ~w5361;
assign w5363 = (pi1007 & ~w5325) | (pi1007 & w10514) | (~w5325 & w10514);
assign w5364 = w5325 & w10515;
assign w5365 = ~w5363 & ~w5364;
assign w5366 = (pi1008 & ~w5062) | (pi1008 & w10516) | (~w5062 & w10516);
assign w5367 = w5062 & w10517;
assign w5368 = ~w5366 & ~w5367;
assign w5369 = (pi1009 & ~w5062) | (pi1009 & w10518) | (~w5062 & w10518);
assign w5370 = w5062 & w10519;
assign w5371 = ~w5369 & ~w5370;
assign w5372 = (pi1010 & ~w5062) | (pi1010 & w10520) | (~w5062 & w10520);
assign w5373 = w5062 & w10521;
assign w5374 = ~w5372 & ~w5373;
assign w5375 = (pi1011 & ~w5062) | (pi1011 & w10522) | (~w5062 & w10522);
assign w5376 = w5062 & w10523;
assign w5377 = ~w5375 & ~w5376;
assign w5378 = w4923 & w10524;
assign w5379 = pi1012 & ~w5378;
assign w5380 = pi2176 & w5378;
assign w5381 = ~w5379 & ~w5380;
assign w5382 = (pi1013 & ~w5062) | (pi1013 & w10525) | (~w5062 & w10525);
assign w5383 = w5062 & w10526;
assign w5384 = ~w5382 & ~w5383;
assign w5385 = ~w5058 & w10527;
assign w5386 = pi1014 & ~w5385;
assign w5387 = pi2189 & w5385;
assign w5388 = ~w5386 & ~w5387;
assign w5389 = (pi1015 & ~w5283) | (pi1015 & w10528) | (~w5283 & w10528);
assign w5390 = w5283 & w10529;
assign w5391 = ~w5389 & ~w5390;
assign w5392 = pi1016 & ~w5385;
assign w5393 = pi2190 & w5385;
assign w5394 = ~w5392 & ~w5393;
assign w5395 = pi1017 & ~w5385;
assign w5396 = pi2182 & w5385;
assign w5397 = ~w5395 & ~w5396;
assign w5398 = ~w5066 & w10530;
assign w5399 = pi1018 & ~w5398;
assign w5400 = pi2196 & w5398;
assign w5401 = ~w5399 & ~w5400;
assign w5402 = ~pi0930 & w5099;
assign w5403 = (pi1019 & ~w5099) | (pi1019 & w10531) | (~w5099 & w10531);
assign w5404 = w5099 & w10532;
assign w5405 = ~w5403 & ~w5404;
assign w5406 = w4930 & w10533;
assign w5407 = pi1020 & ~w5406;
assign w5408 = pi2172 & w5406;
assign w5409 = ~w5407 & ~w5408;
assign w5410 = (pi1021 & ~w5099) | (pi1021 & w10534) | (~w5099 & w10534);
assign w5411 = w5099 & w10433;
assign w5412 = ~w5410 & ~w5411;
assign w5413 = (pi1022 & ~w5099) | (pi1022 & w10535) | (~w5099 & w10535);
assign w5414 = w5099 & w10536;
assign w5415 = ~w5413 & ~w5414;
assign w5416 = (pi1023 & ~w5099) | (pi1023 & w10537) | (~w5099 & w10537);
assign w5417 = w5099 & w10431;
assign w5418 = ~w5416 & ~w5417;
assign w5419 = (pi1024 & ~w5099) | (pi1024 & w10538) | (~w5099 & w10538);
assign w5420 = w5099 & w10539;
assign w5421 = ~w5419 & ~w5420;
assign w5422 = ~pi0941 & w5122;
assign w5423 = (pi1025 & ~w5122) | (pi1025 & w10540) | (~w5122 & w10540);
assign w5424 = w5122 & w10541;
assign w5425 = ~w5423 & ~w5424;
assign w5426 = pi1026 & ~w5385;
assign w5427 = pi2185 & w5385;
assign w5428 = ~w5426 & ~w5427;
assign w5429 = (pi1027 & ~w5066) | (pi1027 & w10542) | (~w5066 & w10542);
assign w5430 = w5066 & w10543;
assign w5431 = ~w5429 & ~w5430;
assign w5432 = (pi1028 & ~w5066) | (pi1028 & w10544) | (~w5066 & w10544);
assign w5433 = w5066 & w10545;
assign w5434 = ~w5432 & ~w5433;
assign w5435 = (pi1029 & ~w5066) | (pi1029 & w10546) | (~w5066 & w10546);
assign w5436 = w5066 & w10547;
assign w5437 = ~w5435 & ~w5436;
assign w5438 = (pi1030 & ~w5325) | (pi1030 & w10548) | (~w5325 & w10548);
assign w5439 = w5325 & w10549;
assign w5440 = ~w5438 & ~w5439;
assign w5441 = (pi1031 & ~w5062) | (pi1031 & w10550) | (~w5062 & w10550);
assign w5442 = w5062 & w10551;
assign w5443 = ~w5441 & ~w5442;
assign w5444 = (pi1032 & ~w5066) | (pi1032 & w10552) | (~w5066 & w10552);
assign w5445 = w5066 & w10553;
assign w5446 = ~w5444 & ~w5445;
assign w5447 = (pi1033 & ~w5066) | (pi1033 & w10554) | (~w5066 & w10554);
assign w5448 = w5066 & w10555;
assign w5449 = ~w5447 & ~w5448;
assign w5450 = (pi1034 & ~w5058) | (pi1034 & w10556) | (~w5058 & w10556);
assign w5451 = w5058 & w10557;
assign w5452 = ~w5450 & ~w5451;
assign w5453 = pi1035 & ~w5406;
assign w5454 = pi2195 & w5406;
assign w5455 = ~w5453 & ~w5454;
assign w5456 = w4930 & w10558;
assign w5457 = pi1036 & ~w5456;
assign w5458 = pi2195 & w5456;
assign w5459 = ~w5457 & ~w5458;
assign w5460 = pi1037 & ~w5385;
assign w5461 = pi2174 & w5385;
assign w5462 = ~w5460 & ~w5461;
assign w5463 = (pi1038 & ~w5122) | (pi1038 & w10559) | (~w5122 & w10559);
assign w5464 = w5122 & w10560;
assign w5465 = ~w5463 & ~w5464;
assign w5466 = pi1039 & ~w5398;
assign w5467 = pi2192 & w5398;
assign w5468 = ~w5466 & ~w5467;
assign w5469 = (pi1040 & ~w5066) | (pi1040 & w10561) | (~w5066 & w10561);
assign w5470 = w5066 & w10562;
assign w5471 = ~w5469 & ~w5470;
assign w5472 = (pi1041 & ~w5066) | (pi1041 & w10563) | (~w5066 & w10563);
assign w5473 = w5066 & w10564;
assign w5474 = ~w5472 & ~w5473;
assign w5475 = pi1042 & ~w5398;
assign w5476 = pi2188 & w5398;
assign w5477 = ~w5475 & ~w5476;
assign w5478 = (pi1043 & ~w5122) | (pi1043 & w10565) | (~w5122 & w10565);
assign w5479 = w5122 & w10489;
assign w5480 = ~w5478 & ~w5479;
assign w5481 = pi1044 & ~w5398;
assign w5482 = pi2177 & w5398;
assign w5483 = ~w5481 & ~w5482;
assign w5484 = pi1045 & ~w5398;
assign w5485 = pi2181 & w5398;
assign w5486 = ~w5484 & ~w5485;
assign w5487 = pi1046 & ~w5398;
assign w5488 = pi2171 & w5398;
assign w5489 = ~w5487 & ~w5488;
assign w5490 = (pi1047 & ~w5283) | (pi1047 & w10566) | (~w5283 & w10566);
assign w5491 = w5283 & w10567;
assign w5492 = ~w5490 & ~w5491;
assign w5493 = pi0941 & w5062;
assign w5494 = (pi1048 & ~w5062) | (pi1048 & w10568) | (~w5062 & w10568);
assign w5495 = w5062 & w10569;
assign w5496 = ~w5494 & ~w5495;
assign w5497 = (pi1049 & ~w5058) | (pi1049 & w10570) | (~w5058 & w10570);
assign w5498 = w5058 & w10571;
assign w5499 = ~w5497 & ~w5498;
assign w5500 = (pi1050 & ~w5122) | (pi1050 & w10572) | (~w5122 & w10572);
assign w5501 = w5122 & w10485;
assign w5502 = ~w5500 & ~w5501;
assign w5503 = (pi1051 & ~w5058) | (pi1051 & w10573) | (~w5058 & w10573);
assign w5504 = w5058 & w10574;
assign w5505 = ~w5503 & ~w5504;
assign w5506 = pi1052 & ~w5398;
assign w5507 = pi2168 & w5398;
assign w5508 = ~w5506 & ~w5507;
assign w5509 = (pi1053 & ~w5066) | (pi1053 & w10575) | (~w5066 & w10575);
assign w5510 = w5066 & w10576;
assign w5511 = ~w5509 & ~w5510;
assign w5512 = (pi1054 & ~w5066) | (pi1054 & w10577) | (~w5066 & w10577);
assign w5513 = w5066 & w10578;
assign w5514 = ~w5512 & ~w5513;
assign w5515 = (pi1055 & ~w5066) | (pi1055 & w10579) | (~w5066 & w10579);
assign w5516 = w5066 & w10580;
assign w5517 = ~w5515 & ~w5516;
assign w5518 = (pi1056 & ~w5066) | (pi1056 & w10581) | (~w5066 & w10581);
assign w5519 = w5066 & w10582;
assign w5520 = ~w5518 & ~w5519;
assign w5521 = (pi1057 & ~w5058) | (pi1057 & w10583) | (~w5058 & w10583);
assign w5522 = w5058 & w10584;
assign w5523 = ~w5521 & ~w5522;
assign w5524 = (pi1058 & ~w5062) | (pi1058 & w10585) | (~w5062 & w10585);
assign w5525 = w5062 & w10586;
assign w5526 = ~w5524 & ~w5525;
assign w5527 = (pi1059 & ~w5058) | (pi1059 & w10587) | (~w5058 & w10587);
assign w5528 = w5058 & w10588;
assign w5529 = ~w5527 & ~w5528;
assign w5530 = (pi1060 & ~w5066) | (pi1060 & w10589) | (~w5066 & w10589);
assign w5531 = w5066 & w10590;
assign w5532 = ~w5530 & ~w5531;
assign w5533 = (pi1061 & ~w5066) | (pi1061 & w10591) | (~w5066 & w10591);
assign w5534 = w5066 & w10592;
assign w5535 = ~w5533 & ~w5534;
assign w5536 = (pi1062 & ~w5283) | (pi1062 & w10593) | (~w5283 & w10593);
assign w5537 = w5283 & w10594;
assign w5538 = ~w5536 & ~w5537;
assign w5539 = (pi1063 & ~w5078) | (pi1063 & w10595) | (~w5078 & w10595);
assign w5540 = w5078 & w10596;
assign w5541 = ~w5539 & ~w5540;
assign w5542 = (pi1064 & ~w5122) | (pi1064 & w10597) | (~w5122 & w10597);
assign w5543 = w5122 & w10598;
assign w5544 = ~w5542 & ~w5543;
assign w5545 = (pi1065 & ~w5066) | (pi1065 & w10599) | (~w5066 & w10599);
assign w5546 = w5066 & w10600;
assign w5547 = ~w5545 & ~w5546;
assign w5548 = (pi1066 & ~w5078) | (pi1066 & w10601) | (~w5078 & w10601);
assign w5549 = w5078 & w10602;
assign w5550 = ~w5548 & ~w5549;
assign w5551 = (pi1067 & ~w5058) | (pi1067 & w10603) | (~w5058 & w10603);
assign w5552 = w5058 & w10604;
assign w5553 = ~w5551 & ~w5552;
assign w5554 = (pi1068 & ~w5058) | (pi1068 & w10605) | (~w5058 & w10605);
assign w5555 = w5058 & w10606;
assign w5556 = ~w5554 & ~w5555;
assign w5557 = (pi1069 & ~w5122) | (pi1069 & w10607) | (~w5122 & w10607);
assign w5558 = w5122 & w10608;
assign w5559 = ~w5557 & ~w5558;
assign w5560 = (pi1070 & ~w5122) | (pi1070 & w10609) | (~w5122 & w10609);
assign w5561 = w5122 & w10610;
assign w5562 = ~w5560 & ~w5561;
assign w5563 = (pi1071 & ~w5122) | (pi1071 & w10611) | (~w5122 & w10611);
assign w5564 = w5122 & w10612;
assign w5565 = ~w5563 & ~w5564;
assign w5566 = (pi1072 & ~w5122) | (pi1072 & w10613) | (~w5122 & w10613);
assign w5567 = w5122 & w10614;
assign w5568 = ~w5566 & ~w5567;
assign w5569 = (pi1073 & ~w5283) | (pi1073 & w10615) | (~w5283 & w10615);
assign w5570 = w5283 & w10616;
assign w5571 = ~w5569 & ~w5570;
assign w5572 = (pi1074 & ~w5122) | (pi1074 & w10617) | (~w5122 & w10617);
assign w5573 = w5122 & w10618;
assign w5574 = ~w5572 & ~w5573;
assign w5575 = (pi1081 & ~w5074) | (pi1081 & w10619) | (~w5074 & w10619);
assign w5576 = w5074 & w10620;
assign w5577 = ~w5575 & ~w5576;
assign w5578 = (pi1082 & ~w5058) | (pi1082 & w10621) | (~w5058 & w10621);
assign w5579 = w5058 & w10622;
assign w5580 = ~w5578 & ~w5579;
assign w5581 = (pi1083 & ~w5078) | (pi1083 & w10623) | (~w5078 & w10623);
assign w5582 = w5078 & w10624;
assign w5583 = ~w5581 & ~w5582;
assign w5584 = (pi1084 & ~w5122) | (pi1084 & w10625) | (~w5122 & w10625);
assign w5585 = w5122 & w10626;
assign w5586 = ~w5584 & ~w5585;
assign w5587 = (pi1085 & ~w5122) | (pi1085 & w10627) | (~w5122 & w10627);
assign w5588 = w5122 & w10628;
assign w5589 = ~w5587 & ~w5588;
assign w5590 = (pi1086 & ~w5062) | (pi1086 & w10629) | (~w5062 & w10629);
assign w5591 = w5062 & w10630;
assign w5592 = ~w5590 & ~w5591;
assign w5593 = (pi1087 & ~w5283) | (pi1087 & w10631) | (~w5283 & w10631);
assign w5594 = w5283 & w10632;
assign w5595 = ~w5593 & ~w5594;
assign w5596 = (pi1088 & ~w5078) | (pi1088 & w10633) | (~w5078 & w10633);
assign w5597 = w5078 & w10634;
assign w5598 = ~w5596 & ~w5597;
assign w5599 = (pi1089 & ~w5078) | (pi1089 & w10635) | (~w5078 & w10635);
assign w5600 = w5078 & w10636;
assign w5601 = ~w5599 & ~w5600;
assign w5602 = (pi1090 & ~w5078) | (pi1090 & w10637) | (~w5078 & w10637);
assign w5603 = w5078 & w10638;
assign w5604 = ~w5602 & ~w5603;
assign w5605 = (pi1091 & ~w5062) | (pi1091 & w10639) | (~w5062 & w10639);
assign w5606 = w5062 & w10640;
assign w5607 = ~w5605 & ~w5606;
assign w5608 = (pi1092 & ~w5062) | (pi1092 & w10641) | (~w5062 & w10641);
assign w5609 = w5062 & w10610;
assign w5610 = ~w5608 & ~w5609;
assign w5611 = (pi1093 & ~w5062) | (pi1093 & w10642) | (~w5062 & w10642);
assign w5612 = w5062 & w10643;
assign w5613 = ~w5611 & ~w5612;
assign w5614 = (pi1094 & ~w5058) | (pi1094 & w10644) | (~w5058 & w10644);
assign w5615 = w5058 & w10645;
assign w5616 = ~w5614 & ~w5615;
assign w5617 = (pi1095 & ~w5058) | (pi1095 & w10646) | (~w5058 & w10646);
assign w5618 = w5058 & w10647;
assign w5619 = ~w5617 & ~w5618;
assign w5620 = (pi1096 & ~w5078) | (pi1096 & w10648) | (~w5078 & w10648);
assign w5621 = w5078 & w10649;
assign w5622 = ~w5620 & ~w5621;
assign w5623 = (pi1097 & ~w5078) | (pi1097 & w10650) | (~w5078 & w10650);
assign w5624 = w5078 & w10651;
assign w5625 = ~w5623 & ~w5624;
assign w5626 = (pi1098 & ~w5058) | (pi1098 & w10652) | (~w5058 & w10652);
assign w5627 = w5058 & w10653;
assign w5628 = ~w5626 & ~w5627;
assign w5629 = (pi1099 & ~w5062) | (pi1099 & w10654) | (~w5062 & w10654);
assign w5630 = w5062 & w10628;
assign w5631 = ~w5629 & ~w5630;
assign w5632 = (pi1100 & ~w5058) | (pi1100 & w10655) | (~w5058 & w10655);
assign w5633 = w5058 & w10656;
assign w5634 = ~w5632 & ~w5633;
assign w5635 = (pi1101 & ~w5283) | (pi1101 & w10657) | (~w5283 & w10657);
assign w5636 = w5283 & w10658;
assign w5637 = ~w5635 & ~w5636;
assign w5638 = (pi1102 & ~w5283) | (pi1102 & w10659) | (~w5283 & w10659);
assign w5639 = w5283 & w10660;
assign w5640 = ~w5638 & ~w5639;
assign w5641 = (pi1103 & ~w5058) | (pi1103 & w10661) | (~w5058 & w10661);
assign w5642 = w5058 & w10662;
assign w5643 = ~w5641 & ~w5642;
assign w5644 = (pi1104 & ~w5058) | (pi1104 & w10663) | (~w5058 & w10663);
assign w5645 = w5058 & w10664;
assign w5646 = ~w5644 & ~w5645;
assign w5647 = ~w5078 & w10665;
assign w5648 = pi1105 & ~w5647;
assign w5649 = pi2190 & w5647;
assign w5650 = ~w5648 & ~w5649;
assign w5651 = pi1106 & ~w5647;
assign w5652 = pi2166 & w5647;
assign w5653 = ~w5651 & ~w5652;
assign w5654 = (pi1107 & ~w5078) | (pi1107 & w10666) | (~w5078 & w10666);
assign w5655 = w5078 & w10667;
assign w5656 = ~w5654 & ~w5655;
assign w5657 = (pi1108 & ~w5058) | (pi1108 & w10668) | (~w5058 & w10668);
assign w5658 = w5058 & w10669;
assign w5659 = ~w5657 & ~w5658;
assign w5660 = (pi1109 & ~w5122) | (pi1109 & w10670) | (~w5122 & w10670);
assign w5661 = w5122 & w10671;
assign w5662 = ~w5660 & ~w5661;
assign w5663 = (pi1110 & ~w5058) | (pi1110 & w10672) | (~w5058 & w10672);
assign w5664 = w5058 & w10673;
assign w5665 = ~w5663 & ~w5664;
assign w5666 = (pi1111 & ~w5058) | (pi1111 & w10674) | (~w5058 & w10674);
assign w5667 = w5058 & w10675;
assign w5668 = ~w5666 & ~w5667;
assign w5669 = pi1112 & ~w5647;
assign w5670 = pi2194 & w5647;
assign w5671 = ~w5669 & ~w5670;
assign w5672 = pi1113 & ~w5647;
assign w5673 = pi2175 & w5647;
assign w5674 = ~w5672 & ~w5673;
assign w5675 = (pi1114 & ~w5122) | (pi1114 & w10676) | (~w5122 & w10676);
assign w5676 = w5122 & w10517;
assign w5677 = ~w5675 & ~w5676;
assign w5678 = pi1115 & ~w5647;
assign w5679 = pi2187 & w5647;
assign w5680 = ~w5678 & ~w5679;
assign w5681 = pi1116 & ~w5647;
assign w5682 = pi2189 & w5647;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = (pi1117 & ~w5074) | (pi1117 & w10677) | (~w5074 & w10677);
assign w5685 = w5074 & w10678;
assign w5686 = ~w5684 & ~w5685;
assign w5687 = (pi1118 & ~w5074) | (pi1118 & w10679) | (~w5074 & w10679);
assign w5688 = w5074 & w10680;
assign w5689 = ~w5687 & ~w5688;
assign w5690 = pi1119 & ~w5647;
assign w5691 = pi2197 & w5647;
assign w5692 = ~w5690 & ~w5691;
assign w5693 = pi1120 & ~w5647;
assign w5694 = pi2183 & w5647;
assign w5695 = ~w5693 & ~w5694;
assign w5696 = pi1121 & ~w5385;
assign w5697 = pi2184 & w5385;
assign w5698 = ~w5696 & ~w5697;
assign w5699 = (pi1122 & ~w5074) | (pi1122 & w10681) | (~w5074 & w10681);
assign w5700 = w5074 & w10682;
assign w5701 = ~w5699 & ~w5700;
assign w5702 = (pi1123 & ~w5078) | (pi1123 & w10683) | (~w5078 & w10683);
assign w5703 = w5078 & w10684;
assign w5704 = ~w5702 & ~w5703;
assign w5705 = (pi1124 & ~w5104) | (pi1124 & w10685) | (~w5104 & w10685);
assign w5706 = w5104 & w10686;
assign w5707 = ~w5705 & ~w5706;
assign w5708 = pi1125 & ~w5378;
assign w5709 = ~pi2194 & w5378;
assign w5710 = ~w5708 & ~w5709;
assign w5711 = pi1126 & ~w5378;
assign w5712 = ~pi2192 & w5378;
assign w5713 = ~w5711 & ~w5712;
assign w5714 = (pi1127 & ~w5078) | (pi1127 & w10687) | (~w5078 & w10687);
assign w5715 = w5078 & w10688;
assign w5716 = ~w5714 & ~w5715;
assign w5717 = pi1128 & ~w5456;
assign w5718 = pi2176 & w5456;
assign w5719 = ~w5717 & ~w5718;
assign w5720 = pi1129 & ~w5378;
assign w5721 = ~pi2197 & w5378;
assign w5722 = ~w5720 & ~w5721;
assign w5723 = pi1130 & ~w5406;
assign w5724 = pi2191 & w5406;
assign w5725 = ~w5723 & ~w5724;
assign w5726 = pi1131 & ~w5406;
assign w5727 = pi2167 & w5406;
assign w5728 = ~w5726 & ~w5727;
assign w5729 = w4914 & w10533;
assign w5730 = pi1132 & ~w5729;
assign w5731 = pi2166 & w5729;
assign w5732 = ~w5730 & ~w5731;
assign w5733 = pi1133 & ~w5729;
assign w5734 = pi2176 & w5729;
assign w5735 = ~w5733 & ~w5734;
assign w5736 = pi1134 & ~w5456;
assign w5737 = pi2172 & w5456;
assign w5738 = ~w5736 & ~w5737;
assign w5739 = (pi1135 & ~w5078) | (pi1135 & w10689) | (~w5078 & w10689);
assign w5740 = w5078 & w10690;
assign w5741 = ~w5739 & ~w5740;
assign w5742 = (pi1136 & ~w5074) | (pi1136 & w10691) | (~w5074 & w10691);
assign w5743 = w5074 & w10692;
assign w5744 = ~w5742 & ~w5743;
assign w5745 = pi1137 & ~w5456;
assign w5746 = pi2178 & w5456;
assign w5747 = ~w5745 & ~w5746;
assign w5748 = pi1138 & ~w5456;
assign w5749 = pi2179 & w5456;
assign w5750 = ~w5748 & ~w5749;
assign w5751 = pi1139 & ~w5378;
assign w5752 = pi2196 & w5378;
assign w5753 = ~w5751 & ~w5752;
assign w5754 = pi1140 & ~w5378;
assign w5755 = pi2193 & w5378;
assign w5756 = ~w5754 & ~w5755;
assign w5757 = pi1141 & ~w5378;
assign w5758 = pi2179 & w5378;
assign w5759 = ~w5757 & ~w5758;
assign w5760 = pi1142 & ~w5378;
assign w5761 = pi2185 & w5378;
assign w5762 = ~w5760 & ~w5761;
assign w5763 = pi1143 & ~w5378;
assign w5764 = pi2187 & w5378;
assign w5765 = ~w5763 & ~w5764;
assign w5766 = pi1144 & ~w5378;
assign w5767 = pi2173 & w5378;
assign w5768 = ~w5766 & ~w5767;
assign w5769 = pi1145 & ~w5456;
assign w5770 = pi2186 & w5456;
assign w5771 = ~w5769 & ~w5770;
assign w5772 = pi1146 & ~w5456;
assign w5773 = pi2183 & w5456;
assign w5774 = ~w5772 & ~w5773;
assign w5775 = pi1147 & ~w5456;
assign w5776 = pi2168 & w5456;
assign w5777 = ~w5775 & ~w5776;
assign w5778 = pi1148 & ~w5456;
assign w5779 = pi2174 & w5456;
assign w5780 = ~w5778 & ~w5779;
assign w5781 = pi1149 & ~w5456;
assign w5782 = pi2197 & w5456;
assign w5783 = ~w5781 & ~w5782;
assign w5784 = pi1150 & ~w5456;
assign w5785 = pi2196 & w5456;
assign w5786 = ~w5784 & ~w5785;
assign w5787 = pi1151 & ~w5456;
assign w5788 = pi2193 & w5456;
assign w5789 = ~w5787 & ~w5788;
assign w5790 = pi1152 & ~w5456;
assign w5791 = pi2189 & w5456;
assign w5792 = ~w5790 & ~w5791;
assign w5793 = pi1153 & ~w5456;
assign w5794 = pi2198 & w5456;
assign w5795 = ~w5793 & ~w5794;
assign w5796 = pi1154 & ~w5456;
assign w5797 = pi2185 & w5456;
assign w5798 = ~w5796 & ~w5797;
assign w5799 = pi1155 & ~w5456;
assign w5800 = pi2187 & w5456;
assign w5801 = ~w5799 & ~w5800;
assign w5802 = pi1156 & ~w5456;
assign w5803 = pi2171 & w5456;
assign w5804 = ~w5802 & ~w5803;
assign w5805 = pi1157 & ~w5456;
assign w5806 = pi2191 & w5456;
assign w5807 = ~w5805 & ~w5806;
assign w5808 = pi1158 & ~w5456;
assign w5809 = pi2194 & w5456;
assign w5810 = ~w5808 & ~w5809;
assign w5811 = pi1159 & ~w5456;
assign w5812 = pi2167 & w5456;
assign w5813 = ~w5811 & ~w5812;
assign w5814 = pi1160 & ~w5456;
assign w5815 = pi2188 & w5456;
assign w5816 = ~w5814 & ~w5815;
assign w5817 = pi1161 & ~w5456;
assign w5818 = pi2184 & w5456;
assign w5819 = ~w5817 & ~w5818;
assign w5820 = pi1162 & ~w5456;
assign w5821 = pi2166 & w5456;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = pi1163 & ~w5456;
assign w5824 = pi2192 & w5456;
assign w5825 = ~w5823 & ~w5824;
assign w5826 = pi1164 & ~w5406;
assign w5827 = pi2186 & w5406;
assign w5828 = ~w5826 & ~w5827;
assign w5829 = pi1165 & ~w5406;
assign w5830 = pi2183 & w5406;
assign w5831 = ~w5829 & ~w5830;
assign w5832 = pi1166 & ~w5406;
assign w5833 = pi2168 & w5406;
assign w5834 = ~w5832 & ~w5833;
assign w5835 = pi1167 & ~w5406;
assign w5836 = pi2174 & w5406;
assign w5837 = ~w5835 & ~w5836;
assign w5838 = pi1168 & ~w5406;
assign w5839 = pi2197 & w5406;
assign w5840 = ~w5838 & ~w5839;
assign w5841 = pi1169 & ~w5406;
assign w5842 = pi2196 & w5406;
assign w5843 = ~w5841 & ~w5842;
assign w5844 = pi1170 & ~w5406;
assign w5845 = pi2193 & w5406;
assign w5846 = ~w5844 & ~w5845;
assign w5847 = pi1171 & ~w5406;
assign w5848 = pi2189 & w5406;
assign w5849 = ~w5847 & ~w5848;
assign w5850 = pi1172 & ~w5406;
assign w5851 = pi2198 & w5406;
assign w5852 = ~w5850 & ~w5851;
assign w5853 = pi1173 & ~w5406;
assign w5854 = pi2185 & w5406;
assign w5855 = ~w5853 & ~w5854;
assign w5856 = pi1174 & ~w5406;
assign w5857 = pi2187 & w5406;
assign w5858 = ~w5856 & ~w5857;
assign w5859 = pi1175 & ~w5406;
assign w5860 = pi2171 & w5406;
assign w5861 = ~w5859 & ~w5860;
assign w5862 = pi1176 & ~w5406;
assign w5863 = pi2169 & w5406;
assign w5864 = ~w5862 & ~w5863;
assign w5865 = pi1177 & ~w5406;
assign w5866 = pi2190 & w5406;
assign w5867 = ~w5865 & ~w5866;
assign w5868 = pi1178 & ~w5406;
assign w5869 = pi2181 & w5406;
assign w5870 = ~w5868 & ~w5869;
assign w5871 = pi1179 & ~w5406;
assign w5872 = pi2182 & w5406;
assign w5873 = ~w5871 & ~w5872;
assign w5874 = pi1180 & ~w5406;
assign w5875 = pi2175 & w5406;
assign w5876 = ~w5874 & ~w5875;
assign w5877 = pi1181 & ~w5406;
assign w5878 = pi2177 & w5406;
assign w5879 = ~w5877 & ~w5878;
assign w5880 = pi1182 & ~w5406;
assign w5881 = pi2173 & w5406;
assign w5882 = ~w5880 & ~w5881;
assign w5883 = pi1183 & ~w5406;
assign w5884 = pi2194 & w5406;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = pi1184 & ~w5406;
assign w5887 = pi2188 & w5406;
assign w5888 = ~w5886 & ~w5887;
assign w5889 = pi1185 & ~w5406;
assign w5890 = pi2184 & w5406;
assign w5891 = ~w5889 & ~w5890;
assign w5892 = pi1186 & ~w5406;
assign w5893 = pi2166 & w5406;
assign w5894 = ~w5892 & ~w5893;
assign w5895 = pi1187 & ~w5406;
assign w5896 = pi2192 & w5406;
assign w5897 = ~w5895 & ~w5896;
assign w5898 = pi1188 & ~w5729;
assign w5899 = pi2186 & w5729;
assign w5900 = ~w5898 & ~w5899;
assign w5901 = pi1189 & ~w5729;
assign w5902 = pi2183 & w5729;
assign w5903 = ~w5901 & ~w5902;
assign w5904 = pi1190 & ~w5729;
assign w5905 = pi2172 & w5729;
assign w5906 = ~w5904 & ~w5905;
assign w5907 = pi1191 & ~w5729;
assign w5908 = pi2168 & w5729;
assign w5909 = ~w5907 & ~w5908;
assign w5910 = pi1192 & ~w5729;
assign w5911 = pi2174 & w5729;
assign w5912 = ~w5910 & ~w5911;
assign w5913 = pi1193 & ~w5729;
assign w5914 = pi2197 & w5729;
assign w5915 = ~w5913 & ~w5914;
assign w5916 = pi1194 & ~w5729;
assign w5917 = pi2196 & w5729;
assign w5918 = ~w5916 & ~w5917;
assign w5919 = pi1195 & ~w5729;
assign w5920 = pi2193 & w5729;
assign w5921 = ~w5919 & ~w5920;
assign w5922 = pi1196 & ~w5729;
assign w5923 = pi2189 & w5729;
assign w5924 = ~w5922 & ~w5923;
assign w5925 = pi1197 & ~w5729;
assign w5926 = pi2179 & w5729;
assign w5927 = ~w5925 & ~w5926;
assign w5928 = pi1198 & ~w5729;
assign w5929 = pi2198 & w5729;
assign w5930 = ~w5928 & ~w5929;
assign w5931 = pi1199 & ~w5729;
assign w5932 = pi2185 & w5729;
assign w5933 = ~w5931 & ~w5932;
assign w5934 = pi1200 & ~w5729;
assign w5935 = pi2187 & w5729;
assign w5936 = ~w5934 & ~w5935;
assign w5937 = pi1201 & ~w5729;
assign w5938 = pi2171 & w5729;
assign w5939 = ~w5937 & ~w5938;
assign w5940 = pi1202 & ~w5729;
assign w5941 = pi2169 & w5729;
assign w5942 = ~w5940 & ~w5941;
assign w5943 = pi1203 & ~w5729;
assign w5944 = pi2190 & w5729;
assign w5945 = ~w5943 & ~w5944;
assign w5946 = pi1204 & ~w5729;
assign w5947 = pi2181 & w5729;
assign w5948 = ~w5946 & ~w5947;
assign w5949 = pi1205 & ~w5729;
assign w5950 = pi2182 & w5729;
assign w5951 = ~w5949 & ~w5950;
assign w5952 = pi1206 & ~w5729;
assign w5953 = pi2191 & w5729;
assign w5954 = ~w5952 & ~w5953;
assign w5955 = pi1207 & ~w5729;
assign w5956 = pi2188 & w5729;
assign w5957 = ~w5955 & ~w5956;
assign w5958 = pi1208 & ~w5729;
assign w5959 = pi2184 & w5729;
assign w5960 = ~w5958 & ~w5959;
assign w5961 = pi1209 & ~w5729;
assign w5962 = pi2192 & w5729;
assign w5963 = ~w5961 & ~w5962;
assign w5964 = pi1210 & ~w5729;
assign w5965 = pi2167 & w5729;
assign w5966 = ~w5964 & ~w5965;
assign w5967 = pi1211 & ~w5729;
assign w5968 = pi2178 & w5729;
assign w5969 = ~w5967 & ~w5968;
assign w5970 = pi1212 & ~w5378;
assign w5971 = ~pi2186 & w5378;
assign w5972 = ~w5970 & ~w5971;
assign w5973 = pi1213 & ~w5378;
assign w5974 = ~pi2183 & w5378;
assign w5975 = ~w5973 & ~w5974;
assign w5976 = pi1214 & ~w5378;
assign w5977 = ~pi2172 & w5378;
assign w5978 = ~w5976 & ~w5977;
assign w5979 = pi1215 & ~w5378;
assign w5980 = ~pi2168 & w5378;
assign w5981 = ~w5979 & ~w5980;
assign w5982 = pi1216 & ~w5378;
assign w5983 = ~pi2174 & w5378;
assign w5984 = ~w5982 & ~w5983;
assign w5985 = pi1217 & ~w5378;
assign w5986 = ~pi2178 & w5378;
assign w5987 = ~w5985 & ~w5986;
assign w5988 = pi1218 & ~w5378;
assign w5989 = ~pi2198 & w5378;
assign w5990 = ~w5988 & ~w5989;
assign w5991 = pi1219 & ~w5378;
assign w5992 = ~pi2191 & w5378;
assign w5993 = ~w5991 & ~w5992;
assign w5994 = pi1220 & ~w5378;
assign w5995 = ~pi2167 & w5378;
assign w5996 = ~w5994 & ~w5995;
assign w5997 = pi1221 & ~w5378;
assign w5998 = ~pi2188 & w5378;
assign w5999 = ~w5997 & ~w5998;
assign w6000 = pi1222 & ~w5378;
assign w6001 = ~pi2184 & w5378;
assign w6002 = ~w6000 & ~w6001;
assign w6003 = pi1223 & ~w5378;
assign w6004 = ~pi2195 & w5378;
assign w6005 = ~w6003 & ~w6004;
assign w6006 = pi1224 & ~w5385;
assign w6007 = pi2167 & w5385;
assign w6008 = ~w6006 & ~w6007;
assign w6009 = (pi1225 & ~w5122) | (pi1225 & w10693) | (~w5122 & w10693);
assign w6010 = w5122 & w10694;
assign w6011 = ~w6009 & ~w6010;
assign w6012 = pi1226 & ~w5385;
assign w6013 = pi2188 & w5385;
assign w6014 = ~w6012 & ~w6013;
assign w6015 = (pi1227 & ~w5122) | (pi1227 & w10695) | (~w5122 & w10695);
assign w6016 = w5122 & w10519;
assign w6017 = ~w6015 & ~w6016;
assign w6018 = pi1228 & ~w5385;
assign w6019 = pi2166 & w5385;
assign w6020 = ~w6018 & ~w6019;
assign w6021 = pi1229 & ~w5385;
assign w6022 = pi2195 & w5385;
assign w6023 = ~w6021 & ~w6022;
assign w6024 = pi1230 & ~w5385;
assign w6025 = pi2192 & w5385;
assign w6026 = ~w6024 & ~w6025;
assign w6027 = (pi1231 & ~w5058) | (pi1231 & w10696) | (~w5058 & w10696);
assign w6028 = w5058 & w10697;
assign w6029 = ~w6027 & ~w6028;
assign w6030 = (pi1232 & ~w5122) | (pi1232 & w10698) | (~w5122 & w10698);
assign w6031 = w5122 & w10699;
assign w6032 = ~w6030 & ~w6031;
assign w6033 = (pi1233 & ~w5058) | (pi1233 & w10700) | (~w5058 & w10700);
assign w6034 = w5058 & w10701;
assign w6035 = ~w6033 & ~w6034;
assign w6036 = (pi1234 & ~w5122) | (pi1234 & w10702) | (~w5122 & w10702);
assign w6037 = w5122 & w10703;
assign w6038 = ~w6036 & ~w6037;
assign w6039 = (pi1235 & ~w5058) | (pi1235 & w10704) | (~w5058 & w10704);
assign w6040 = w5058 & w10705;
assign w6041 = ~w6039 & ~w6040;
assign w6042 = (pi1236 & ~w5058) | (pi1236 & w10706) | (~w5058 & w10706);
assign w6043 = w5058 & w10707;
assign w6044 = ~w6042 & ~w6043;
assign w6045 = (pi1237 & ~w5122) | (pi1237 & w10708) | (~w5122 & w10708);
assign w6046 = w5122 & w10709;
assign w6047 = ~w6045 & ~w6046;
assign w6048 = (pi1238 & ~w5058) | (pi1238 & w10710) | (~w5058 & w10710);
assign w6049 = w5058 & w10711;
assign w6050 = ~w6048 & ~w6049;
assign w6051 = (pi1239 & ~w5058) | (pi1239 & w10712) | (~w5058 & w10712);
assign w6052 = w5058 & w10713;
assign w6053 = ~w6051 & ~w6052;
assign w6054 = (pi1240 & ~w5058) | (pi1240 & w10714) | (~w5058 & w10714);
assign w6055 = w5058 & w10715;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = (pi1241 & ~w5122) | (pi1241 & w10716) | (~w5122 & w10716);
assign w6058 = w5122 & w10523;
assign w6059 = ~w6057 & ~w6058;
assign w6060 = (pi1242 & ~w5058) | (pi1242 & w10717) | (~w5058 & w10717);
assign w6061 = w5058 & w10718;
assign w6062 = ~w6060 & ~w6061;
assign w6063 = (pi1243 & ~w5122) | (pi1243 & w10719) | (~w5122 & w10719);
assign w6064 = w5122 & w10521;
assign w6065 = ~w6063 & ~w6064;
assign w6066 = (pi1244 & ~w5058) | (pi1244 & w10720) | (~w5058 & w10720);
assign w6067 = w5058 & w10721;
assign w6068 = ~w6066 & ~w6067;
assign w6069 = (pi1245 & ~w5122) | (pi1245 & w10722) | (~w5122 & w10722);
assign w6070 = w5122 & w10723;
assign w6071 = ~w6069 & ~w6070;
assign w6072 = (pi1246 & ~w5058) | (pi1246 & w10724) | (~w5058 & w10724);
assign w6073 = w5058 & w10725;
assign w6074 = ~w6072 & ~w6073;
assign w6075 = (pi1247 & ~w5058) | (pi1247 & w10726) | (~w5058 & w10726);
assign w6076 = w5058 & w10727;
assign w6077 = ~w6075 & ~w6076;
assign w6078 = (pi1248 & ~w5122) | (pi1248 & w10728) | (~w5122 & w10728);
assign w6079 = w5122 & w10729;
assign w6080 = ~w6078 & ~w6079;
assign w6081 = (pi1249 & ~w5058) | (pi1249 & w10730) | (~w5058 & w10730);
assign w6082 = w5058 & w10731;
assign w6083 = ~w6081 & ~w6082;
assign w6084 = (pi1250 & ~w5058) | (pi1250 & w10732) | (~w5058 & w10732);
assign w6085 = w5058 & w10733;
assign w6086 = ~w6084 & ~w6085;
assign w6087 = (pi1251 & ~w5122) | (pi1251 & w10734) | (~w5122 & w10734);
assign w6088 = w5122 & w10735;
assign w6089 = ~w6087 & ~w6088;
assign w6090 = (pi1252 & ~w5058) | (pi1252 & w10736) | (~w5058 & w10736);
assign w6091 = w5058 & w10737;
assign w6092 = ~w6090 & ~w6091;
assign w6093 = (pi1253 & ~w5062) | (pi1253 & w10738) | (~w5062 & w10738);
assign w6094 = w5062 & w10739;
assign w6095 = ~w6093 & ~w6094;
assign w6096 = (pi1254 & ~w5058) | (pi1254 & w10740) | (~w5058 & w10740);
assign w6097 = pi2181 & w5117;
assign w6098 = ~w6096 & ~w6097;
assign w6099 = pi1255 & ~w5493;
assign w6100 = pi2183 & w5493;
assign w6101 = ~w6099 & ~w6100;
assign w6102 = pi1256 & ~w5117;
assign w6103 = pi2175 & w5117;
assign w6104 = ~w6102 & ~w6103;
assign w6105 = pi1257 & ~w5117;
assign w6106 = pi2191 & w5117;
assign w6107 = ~w6105 & ~w6106;
assign w6108 = pi1258 & ~w5117;
assign w6109 = pi2177 & w5117;
assign w6110 = ~w6108 & ~w6109;
assign w6111 = pi1259 & ~w5117;
assign w6112 = pi2173 & w5117;
assign w6113 = ~w6111 & ~w6112;
assign w6114 = pi1260 & ~w5493;
assign w6115 = pi2168 & w5493;
assign w6116 = ~w6114 & ~w6115;
assign w6117 = pi1261 & ~w5117;
assign w6118 = pi2167 & w5117;
assign w6119 = ~w6117 & ~w6118;
assign w6120 = pi1262 & ~w5493;
assign w6121 = pi2174 & w5493;
assign w6122 = ~w6120 & ~w6121;
assign w6123 = pi1263 & ~w5117;
assign w6124 = pi2188 & w5117;
assign w6125 = ~w6123 & ~w6124;
assign w6126 = pi1264 & ~w5493;
assign w6127 = pi2197 & w5493;
assign w6128 = ~w6126 & ~w6127;
assign w6129 = pi1265 & ~w5117;
assign w6130 = pi2166 & w5117;
assign w6131 = ~w6129 & ~w6130;
assign w6132 = pi1266 & ~w5493;
assign w6133 = pi2178 & w5493;
assign w6134 = ~w6132 & ~w6133;
assign w6135 = pi1267 & ~w5117;
assign w6136 = pi2192 & w5117;
assign w6137 = ~w6135 & ~w6136;
assign w6138 = pi1268 & ~w5493;
assign w6139 = pi2196 & w5493;
assign w6140 = ~w6138 & ~w6139;
assign w6141 = pi1269 & ~w5493;
assign w6142 = pi2193 & w5493;
assign w6143 = ~w6141 & ~w6142;
assign w6144 = pi1270 & ~w5493;
assign w6145 = pi2179 & w5493;
assign w6146 = ~w6144 & ~w6145;
assign w6147 = pi1271 & ~w5493;
assign w6148 = pi2198 & w5493;
assign w6149 = ~w6147 & ~w6148;
assign w6150 = pi1272 & ~w5493;
assign w6151 = pi2187 & w5493;
assign w6152 = ~w6150 & ~w6151;
assign w6153 = pi1273 & ~w5493;
assign w6154 = pi2171 & w5493;
assign w6155 = ~w6153 & ~w6154;
assign w6156 = pi1274 & ~w5493;
assign w6157 = pi2169 & w5493;
assign w6158 = ~w6156 & ~w6157;
assign w6159 = pi1275 & ~w5493;
assign w6160 = pi2190 & w5493;
assign w6161 = ~w6159 & ~w6160;
assign w6162 = pi1276 & ~w5493;
assign w6163 = pi2181 & w5493;
assign w6164 = ~w6162 & ~w6163;
assign w6165 = pi1277 & ~w5493;
assign w6166 = pi2182 & w5493;
assign w6167 = ~w6165 & ~w6166;
assign w6168 = pi1278 & ~w5493;
assign w6169 = pi2175 & w5493;
assign w6170 = ~w6168 & ~w6169;
assign w6171 = pi1279 & ~w5493;
assign w6172 = pi2177 & w5493;
assign w6173 = ~w6171 & ~w6172;
assign w6174 = pi1280 & ~w5493;
assign w6175 = pi2173 & w5493;
assign w6176 = ~w6174 & ~w6175;
assign w6177 = pi1281 & ~w5493;
assign w6178 = pi2194 & w5493;
assign w6179 = ~w6177 & ~w6178;
assign w6180 = pi1282 & ~w5493;
assign w6181 = pi2167 & w5493;
assign w6182 = ~w6180 & ~w6181;
assign w6183 = pi1283 & ~w5493;
assign w6184 = pi2188 & w5493;
assign w6185 = ~w6183 & ~w6184;
assign w6186 = pi1284 & ~w5493;
assign w6187 = pi2184 & w5493;
assign w6188 = ~w6186 & ~w6187;
assign w6189 = pi1285 & ~w5493;
assign w6190 = pi2166 & w5493;
assign w6191 = ~w6189 & ~w6190;
assign w6192 = pi1286 & ~w5493;
assign w6193 = pi2192 & w5493;
assign w6194 = ~w6192 & ~w6193;
assign w6195 = pi1287 & ~w5123;
assign w6196 = pi2186 & w5123;
assign w6197 = ~w6195 & ~w6196;
assign w6198 = pi1288 & ~w5123;
assign w6199 = pi2183 & w5123;
assign w6200 = ~w6198 & ~w6199;
assign w6201 = pi1289 & ~w5123;
assign w6202 = pi2168 & w5123;
assign w6203 = ~w6201 & ~w6202;
assign w6204 = pi1290 & ~w5123;
assign w6205 = pi2174 & w5123;
assign w6206 = ~w6204 & ~w6205;
assign w6207 = pi1291 & ~w5123;
assign w6208 = pi2197 & w5123;
assign w6209 = ~w6207 & ~w6208;
assign w6210 = pi1292 & ~w5123;
assign w6211 = pi2196 & w5123;
assign w6212 = ~w6210 & ~w6211;
assign w6213 = pi1293 & ~w5123;
assign w6214 = pi2193 & w5123;
assign w6215 = ~w6213 & ~w6214;
assign w6216 = pi1294 & ~w5123;
assign w6217 = pi2189 & w5123;
assign w6218 = ~w6216 & ~w6217;
assign w6219 = pi1295 & ~w5123;
assign w6220 = pi2198 & w5123;
assign w6221 = ~w6219 & ~w6220;
assign w6222 = pi1296 & ~w5123;
assign w6223 = pi2185 & w5123;
assign w6224 = ~w6222 & ~w6223;
assign w6225 = pi1297 & ~w5123;
assign w6226 = pi2187 & w5123;
assign w6227 = ~w6225 & ~w6226;
assign w6228 = pi1298 & ~w5123;
assign w6229 = pi2171 & w5123;
assign w6230 = ~w6228 & ~w6229;
assign w6231 = pi1299 & ~w5123;
assign w6232 = pi2169 & w5123;
assign w6233 = ~w6231 & ~w6232;
assign w6234 = pi1300 & ~w5123;
assign w6235 = pi2170 & w5123;
assign w6236 = ~w6234 & ~w6235;
assign w6237 = pi1301 & ~w5123;
assign w6238 = pi2182 & w5123;
assign w6239 = ~w6237 & ~w6238;
assign w6240 = pi1302 & ~w5123;
assign w6241 = pi2175 & w5123;
assign w6242 = ~w6240 & ~w6241;
assign w6243 = pi1303 & ~w5123;
assign w6244 = pi2191 & w5123;
assign w6245 = ~w6243 & ~w6244;
assign w6246 = pi1304 & ~w5123;
assign w6247 = pi2173 & w5123;
assign w6248 = ~w6246 & ~w6247;
assign w6249 = pi1305 & ~w5123;
assign w6250 = pi2167 & w5123;
assign w6251 = ~w6249 & ~w6250;
assign w6252 = pi1306 & ~w5123;
assign w6253 = pi2188 & w5123;
assign w6254 = ~w6252 & ~w6253;
assign w6255 = pi1307 & ~w5123;
assign w6256 = pi2166 & w5123;
assign w6257 = ~w6255 & ~w6256;
assign w6258 = pi1308 & ~w5123;
assign w6259 = pi2192 & w5123;
assign w6260 = ~w6258 & ~w6259;
assign w6261 = pi1309 & ~w5123;
assign w6262 = pi2190 & w5123;
assign w6263 = ~w6261 & ~w6262;
assign w6264 = pi1310 & ~w5159;
assign w6265 = pi2186 & w5159;
assign w6266 = ~w6264 & ~w6265;
assign w6267 = pi1311 & ~w5159;
assign w6268 = pi2183 & w5159;
assign w6269 = ~w6267 & ~w6268;
assign w6270 = pi1312 & ~w5159;
assign w6271 = pi2172 & w5159;
assign w6272 = ~w6270 & ~w6271;
assign w6273 = pi1313 & ~w5159;
assign w6274 = pi2174 & w5159;
assign w6275 = ~w6273 & ~w6274;
assign w6276 = pi1314 & ~w5159;
assign w6277 = pi2197 & w5159;
assign w6278 = ~w6276 & ~w6277;
assign w6279 = pi1315 & ~w5159;
assign w6280 = pi2178 & w5159;
assign w6281 = ~w6279 & ~w6280;
assign w6282 = pi1316 & ~w5159;
assign w6283 = pi2193 & w5159;
assign w6284 = ~w6282 & ~w6283;
assign w6285 = pi1317 & ~w5159;
assign w6286 = pi2189 & w5159;
assign w6287 = ~w6285 & ~w6286;
assign w6288 = pi1318 & ~w5159;
assign w6289 = pi2179 & w5159;
assign w6290 = ~w6288 & ~w6289;
assign w6291 = pi1319 & ~w5159;
assign w6292 = pi2198 & w5159;
assign w6293 = ~w6291 & ~w6292;
assign w6294 = pi1320 & ~w5159;
assign w6295 = pi2185 & w5159;
assign w6296 = ~w6294 & ~w6295;
assign w6297 = pi1321 & ~w5159;
assign w6298 = pi2187 & w5159;
assign w6299 = ~w6297 & ~w6298;
assign w6300 = pi1322 & ~w5159;
assign w6301 = pi2176 & w5159;
assign w6302 = ~w6300 & ~w6301;
assign w6303 = pi1323 & ~w5159;
assign w6304 = pi2169 & w5159;
assign w6305 = ~w6303 & ~w6304;
assign w6306 = pi1324 & ~w5159;
assign w6307 = pi2190 & w5159;
assign w6308 = ~w6306 & ~w6307;
assign w6309 = pi1325 & ~w5159;
assign w6310 = pi2170 & w5159;
assign w6311 = ~w6309 & ~w6310;
assign w6312 = pi1326 & ~w5159;
assign w6313 = pi2182 & w5159;
assign w6314 = ~w6312 & ~w6313;
assign w6315 = pi1327 & ~w5159;
assign w6316 = pi2175 & w5159;
assign w6317 = ~w6315 & ~w6316;
assign w6318 = pi1328 & ~w5159;
assign w6319 = pi2191 & w5159;
assign w6320 = ~w6318 & ~w6319;
assign w6321 = pi1329 & ~w5159;
assign w6322 = pi2173 & w5159;
assign w6323 = ~w6321 & ~w6322;
assign w6324 = pi1330 & ~w5159;
assign w6325 = pi2194 & w5159;
assign w6326 = ~w6324 & ~w6325;
assign w6327 = pi1331 & ~w5159;
assign w6328 = pi2167 & w5159;
assign w6329 = ~w6327 & ~w6328;
assign w6330 = pi1332 & ~w5159;
assign w6331 = pi2184 & w5159;
assign w6332 = ~w6330 & ~w6331;
assign w6333 = pi1333 & ~w5159;
assign w6334 = pi2166 & w5159;
assign w6335 = ~w6333 & ~w6334;
assign w6336 = pi1334 & ~w5159;
assign w6337 = pi2195 & w5159;
assign w6338 = ~w6336 & ~w6337;
assign w6339 = pi1335 & ~w5398;
assign w6340 = pi2186 & w5398;
assign w6341 = ~w6339 & ~w6340;
assign w6342 = pi1336 & ~w5398;
assign w6343 = pi2183 & w5398;
assign w6344 = ~w6342 & ~w6343;
assign w6345 = pi1337 & ~w5398;
assign w6346 = pi2172 & w5398;
assign w6347 = ~w6345 & ~w6346;
assign w6348 = pi1338 & ~w5398;
assign w6349 = pi2174 & w5398;
assign w6350 = ~w6348 & ~w6349;
assign w6351 = pi1339 & ~w5398;
assign w6352 = pi2197 & w5398;
assign w6353 = ~w6351 & ~w6352;
assign w6354 = pi1340 & ~w5398;
assign w6355 = pi2178 & w5398;
assign w6356 = ~w6354 & ~w6355;
assign w6357 = pi1341 & ~w5398;
assign w6358 = pi2193 & w5398;
assign w6359 = ~w6357 & ~w6358;
assign w6360 = pi1342 & ~w5398;
assign w6361 = pi2189 & w5398;
assign w6362 = ~w6360 & ~w6361;
assign w6363 = pi1343 & ~w5398;
assign w6364 = pi2179 & w5398;
assign w6365 = ~w6363 & ~w6364;
assign w6366 = pi1344 & ~w5398;
assign w6367 = pi2198 & w5398;
assign w6368 = ~w6366 & ~w6367;
assign w6369 = pi1345 & ~w5398;
assign w6370 = pi2185 & w5398;
assign w6371 = ~w6369 & ~w6370;
assign w6372 = pi1346 & ~w5398;
assign w6373 = pi2187 & w5398;
assign w6374 = ~w6372 & ~w6373;
assign w6375 = pi1347 & ~w5398;
assign w6376 = pi2176 & w5398;
assign w6377 = ~w6375 & ~w6376;
assign w6378 = pi1348 & ~w5398;
assign w6379 = pi2169 & w5398;
assign w6380 = ~w6378 & ~w6379;
assign w6381 = pi1349 & ~w5398;
assign w6382 = pi2190 & w5398;
assign w6383 = ~w6381 & ~w6382;
assign w6384 = pi1350 & ~w5398;
assign w6385 = pi2170 & w5398;
assign w6386 = ~w6384 & ~w6385;
assign w6387 = pi1351 & ~w5398;
assign w6388 = pi2182 & w5398;
assign w6389 = ~w6387 & ~w6388;
assign w6390 = pi1352 & ~w5398;
assign w6391 = pi2175 & w5398;
assign w6392 = ~w6390 & ~w6391;
assign w6393 = pi1353 & ~w5398;
assign w6394 = pi2191 & w5398;
assign w6395 = ~w6393 & ~w6394;
assign w6396 = pi1354 & ~w5398;
assign w6397 = pi2173 & w5398;
assign w6398 = ~w6396 & ~w6397;
assign w6399 = pi1355 & ~w5398;
assign w6400 = pi2194 & w5398;
assign w6401 = ~w6399 & ~w6400;
assign w6402 = pi1356 & ~w5398;
assign w6403 = pi2167 & w5398;
assign w6404 = ~w6402 & ~w6403;
assign w6405 = pi1357 & ~w5398;
assign w6406 = pi2184 & w5398;
assign w6407 = ~w6405 & ~w6406;
assign w6408 = pi1358 & ~w5398;
assign w6409 = pi2166 & w5398;
assign w6410 = ~w6408 & ~w6409;
assign w6411 = pi1359 & ~w5398;
assign w6412 = pi2195 & w5398;
assign w6413 = ~w6411 & ~w6412;
assign w6414 = pi1360 & ~w5169;
assign w6415 = pi2186 & w5169;
assign w6416 = ~w6414 & ~w6415;
assign w6417 = pi1361 & ~w5169;
assign w6418 = pi2183 & w5169;
assign w6419 = ~w6417 & ~w6418;
assign w6420 = pi1362 & ~w5169;
assign w6421 = pi2172 & w5169;
assign w6422 = ~w6420 & ~w6421;
assign w6423 = pi1363 & ~w5169;
assign w6424 = pi2174 & w5169;
assign w6425 = ~w6423 & ~w6424;
assign w6426 = pi1364 & ~w5169;
assign w6427 = pi2197 & w5169;
assign w6428 = ~w6426 & ~w6427;
assign w6429 = pi1365 & ~w5169;
assign w6430 = pi2178 & w5169;
assign w6431 = ~w6429 & ~w6430;
assign w6432 = pi1366 & ~w5169;
assign w6433 = pi2193 & w5169;
assign w6434 = ~w6432 & ~w6433;
assign w6435 = pi1367 & ~w5169;
assign w6436 = pi2189 & w5169;
assign w6437 = ~w6435 & ~w6436;
assign w6438 = pi1368 & ~w5169;
assign w6439 = pi2179 & w5169;
assign w6440 = ~w6438 & ~w6439;
assign w6441 = pi1369 & ~w5169;
assign w6442 = pi2198 & w5169;
assign w6443 = ~w6441 & ~w6442;
assign w6444 = pi1370 & ~w5169;
assign w6445 = pi2185 & w5169;
assign w6446 = ~w6444 & ~w6445;
assign w6447 = pi1371 & ~w5169;
assign w6448 = pi2187 & w5169;
assign w6449 = ~w6447 & ~w6448;
assign w6450 = pi1372 & ~w5169;
assign w6451 = pi2176 & w5169;
assign w6452 = ~w6450 & ~w6451;
assign w6453 = pi1373 & ~w5169;
assign w6454 = pi2169 & w5169;
assign w6455 = ~w6453 & ~w6454;
assign w6456 = pi1374 & ~w5169;
assign w6457 = pi2190 & w5169;
assign w6458 = ~w6456 & ~w6457;
assign w6459 = pi1375 & ~w5169;
assign w6460 = pi2170 & w5169;
assign w6461 = ~w6459 & ~w6460;
assign w6462 = pi1376 & ~w5169;
assign w6463 = pi2182 & w5169;
assign w6464 = ~w6462 & ~w6463;
assign w6465 = pi1377 & ~w5169;
assign w6466 = pi2175 & w5169;
assign w6467 = ~w6465 & ~w6466;
assign w6468 = pi1378 & ~w5169;
assign w6469 = pi2191 & w5169;
assign w6470 = ~w6468 & ~w6469;
assign w6471 = pi1379 & ~w5169;
assign w6472 = pi2173 & w5169;
assign w6473 = ~w6471 & ~w6472;
assign w6474 = pi1380 & ~w5169;
assign w6475 = pi2194 & w5169;
assign w6476 = ~w6474 & ~w6475;
assign w6477 = pi1381 & ~w5169;
assign w6478 = pi2167 & w5169;
assign w6479 = ~w6477 & ~w6478;
assign w6480 = pi1382 & ~w5169;
assign w6481 = pi2184 & w5169;
assign w6482 = ~w6480 & ~w6481;
assign w6483 = pi1383 & ~w5169;
assign w6484 = pi2166 & w5169;
assign w6485 = ~w6483 & ~w6484;
assign w6486 = pi1384 & ~w5169;
assign w6487 = pi2195 & w5169;
assign w6488 = ~w6486 & ~w6487;
assign w6489 = pi1385 & ~w5493;
assign w6490 = pi2185 & w5493;
assign w6491 = ~w6489 & ~w6490;
assign w6492 = pi1386 & ~w5402;
assign w6493 = pi2186 & w5402;
assign w6494 = ~w6492 & ~w6493;
assign w6495 = pi1387 & ~w5402;
assign w6496 = pi2183 & w5402;
assign w6497 = ~w6495 & ~w6496;
assign w6498 = pi1388 & ~w5402;
assign w6499 = pi2168 & w5402;
assign w6500 = ~w6498 & ~w6499;
assign w6501 = pi1389 & ~w5402;
assign w6502 = pi2174 & w5402;
assign w6503 = ~w6501 & ~w6502;
assign w6504 = pi1390 & ~w5402;
assign w6505 = pi2197 & w5402;
assign w6506 = ~w6504 & ~w6505;
assign w6507 = pi1391 & ~w5166;
assign w6508 = pi2197 & w5166;
assign w6509 = ~w6507 & ~w6508;
assign w6510 = pi1392 & ~w5402;
assign w6511 = pi2196 & w5402;
assign w6512 = ~w6510 & ~w6511;
assign w6513 = pi1393 & ~w5402;
assign w6514 = pi2193 & w5402;
assign w6515 = ~w6513 & ~w6514;
assign w6516 = pi1394 & ~w5402;
assign w6517 = pi2189 & w5402;
assign w6518 = ~w6516 & ~w6517;
assign w6519 = pi1395 & ~w5402;
assign w6520 = pi2198 & w5402;
assign w6521 = ~w6519 & ~w6520;
assign w6522 = pi1396 & ~w5402;
assign w6523 = pi2185 & w5402;
assign w6524 = ~w6522 & ~w6523;
assign w6525 = pi1397 & ~w5402;
assign w6526 = pi2187 & w5402;
assign w6527 = ~w6525 & ~w6526;
assign w6528 = pi1398 & ~w5402;
assign w6529 = pi2171 & w5402;
assign w6530 = ~w6528 & ~w6529;
assign w6531 = pi1399 & ~w5402;
assign w6532 = pi2169 & w5402;
assign w6533 = ~w6531 & ~w6532;
assign w6534 = pi1400 & ~w5402;
assign w6535 = pi2190 & w5402;
assign w6536 = ~w6534 & ~w6535;
assign w6537 = pi1401 & ~w5402;
assign w6538 = pi2181 & w5402;
assign w6539 = ~w6537 & ~w6538;
assign w6540 = pi1402 & ~w5402;
assign w6541 = pi2182 & w5402;
assign w6542 = ~w6540 & ~w6541;
assign w6543 = pi1403 & ~w5402;
assign w6544 = pi2175 & w5402;
assign w6545 = ~w6543 & ~w6544;
assign w6546 = pi1404 & ~w5402;
assign w6547 = pi2177 & w5402;
assign w6548 = ~w6546 & ~w6547;
assign w6549 = pi1405 & ~w5402;
assign w6550 = pi2173 & w5402;
assign w6551 = ~w6549 & ~w6550;
assign w6552 = pi1406 & ~w5402;
assign w6553 = pi2194 & w5402;
assign w6554 = ~w6552 & ~w6553;
assign w6555 = pi1407 & ~w5402;
assign w6556 = pi2188 & w5402;
assign w6557 = ~w6555 & ~w6556;
assign w6558 = pi1408 & ~w5402;
assign w6559 = pi2184 & w5402;
assign w6560 = ~w6558 & ~w6559;
assign w6561 = pi1409 & ~w5402;
assign w6562 = pi2166 & w5402;
assign w6563 = ~w6561 & ~w6562;
assign w6564 = pi1410 & ~w5402;
assign w6565 = pi2192 & w5402;
assign w6566 = ~w6564 & ~w6565;
assign w6567 = pi0930 & w5070;
assign w6568 = pi1411 & ~w6567;
assign w6569 = pi2186 & w6567;
assign w6570 = ~w6568 & ~w6569;
assign w6571 = pi1412 & ~w6567;
assign w6572 = pi2183 & w6567;
assign w6573 = ~w6571 & ~w6572;
assign w6574 = pi1413 & ~w6567;
assign w6575 = pi2168 & w6567;
assign w6576 = ~w6574 & ~w6575;
assign w6577 = pi1414 & ~w6567;
assign w6578 = pi2174 & w6567;
assign w6579 = ~w6577 & ~w6578;
assign w6580 = pi1415 & ~w6567;
assign w6581 = pi2197 & w6567;
assign w6582 = ~w6580 & ~w6581;
assign w6583 = pi1416 & ~w6567;
assign w6584 = pi2196 & w6567;
assign w6585 = ~w6583 & ~w6584;
assign w6586 = pi1417 & ~w6567;
assign w6587 = pi2193 & w6567;
assign w6588 = ~w6586 & ~w6587;
assign w6589 = pi1418 & ~w6567;
assign w6590 = pi2189 & w6567;
assign w6591 = ~w6589 & ~w6590;
assign w6592 = pi1419 & ~w6567;
assign w6593 = pi2198 & w6567;
assign w6594 = ~w6592 & ~w6593;
assign w6595 = pi1420 & ~w6567;
assign w6596 = pi2185 & w6567;
assign w6597 = ~w6595 & ~w6596;
assign w6598 = pi1421 & ~w6567;
assign w6599 = pi2187 & w6567;
assign w6600 = ~w6598 & ~w6599;
assign w6601 = pi1422 & ~w6567;
assign w6602 = pi2171 & w6567;
assign w6603 = ~w6601 & ~w6602;
assign w6604 = pi1423 & ~w6567;
assign w6605 = pi2169 & w6567;
assign w6606 = ~w6604 & ~w6605;
assign w6607 = pi1424 & ~w6567;
assign w6608 = pi2190 & w6567;
assign w6609 = ~w6607 & ~w6608;
assign w6610 = pi1425 & ~w6567;
assign w6611 = pi2181 & w6567;
assign w6612 = ~w6610 & ~w6611;
assign w6613 = pi1426 & ~w6567;
assign w6614 = pi2182 & w6567;
assign w6615 = ~w6613 & ~w6614;
assign w6616 = pi1427 & ~w6567;
assign w6617 = pi2175 & w6567;
assign w6618 = ~w6616 & ~w6617;
assign w6619 = pi1428 & ~w6567;
assign w6620 = pi2177 & w6567;
assign w6621 = ~w6619 & ~w6620;
assign w6622 = pi1429 & ~w6567;
assign w6623 = pi2173 & w6567;
assign w6624 = ~w6622 & ~w6623;
assign w6625 = pi1430 & ~w6567;
assign w6626 = pi2194 & w6567;
assign w6627 = ~w6625 & ~w6626;
assign w6628 = pi1431 & ~w6567;
assign w6629 = pi2167 & w6567;
assign w6630 = ~w6628 & ~w6629;
assign w6631 = pi1432 & ~w6567;
assign w6632 = pi2188 & w6567;
assign w6633 = ~w6631 & ~w6632;
assign w6634 = pi1433 & ~w6567;
assign w6635 = pi2184 & w6567;
assign w6636 = ~w6634 & ~w6635;
assign w6637 = pi1434 & ~w6567;
assign w6638 = pi2166 & w6567;
assign w6639 = ~w6637 & ~w6638;
assign w6640 = pi1435 & ~w6567;
assign w6641 = pi2192 & w6567;
assign w6642 = ~w6640 & ~w6641;
assign w6643 = pi1436 & ~w5100;
assign w6644 = pi2186 & w5100;
assign w6645 = ~w6643 & ~w6644;
assign w6646 = pi1437 & ~w5100;
assign w6647 = pi2183 & w5100;
assign w6648 = ~w6646 & ~w6647;
assign w6649 = pi1438 & ~w5100;
assign w6650 = pi2168 & w5100;
assign w6651 = ~w6649 & ~w6650;
assign w6652 = pi1439 & ~w5100;
assign w6653 = pi2174 & w5100;
assign w6654 = ~w6652 & ~w6653;
assign w6655 = pi1440 & ~w5100;
assign w6656 = pi2197 & w5100;
assign w6657 = ~w6655 & ~w6656;
assign w6658 = pi1441 & ~w5100;
assign w6659 = pi2196 & w5100;
assign w6660 = ~w6658 & ~w6659;
assign w6661 = pi1442 & ~w5100;
assign w6662 = pi2193 & w5100;
assign w6663 = ~w6661 & ~w6662;
assign w6664 = pi1443 & ~w5100;
assign w6665 = pi2189 & w5100;
assign w6666 = ~w6664 & ~w6665;
assign w6667 = pi1444 & ~w5100;
assign w6668 = pi2198 & w5100;
assign w6669 = ~w6667 & ~w6668;
assign w6670 = pi1445 & ~w5100;
assign w6671 = pi2185 & w5100;
assign w6672 = ~w6670 & ~w6671;
assign w6673 = pi1446 & ~w5100;
assign w6674 = pi2187 & w5100;
assign w6675 = ~w6673 & ~w6674;
assign w6676 = pi1447 & ~w5252;
assign w6677 = pi2193 & w5252;
assign w6678 = ~w6676 & ~w6677;
assign w6679 = pi1448 & ~w5100;
assign w6680 = pi2171 & w5100;
assign w6681 = ~w6679 & ~w6680;
assign w6682 = pi1449 & ~w5100;
assign w6683 = pi2169 & w5100;
assign w6684 = ~w6682 & ~w6683;
assign w6685 = pi1450 & ~w5100;
assign w6686 = pi2190 & w5100;
assign w6687 = ~w6685 & ~w6686;
assign w6688 = pi1451 & ~w5100;
assign w6689 = pi2181 & w5100;
assign w6690 = ~w6688 & ~w6689;
assign w6691 = pi1452 & ~w5100;
assign w6692 = pi2182 & w5100;
assign w6693 = ~w6691 & ~w6692;
assign w6694 = pi1453 & ~w5100;
assign w6695 = pi2175 & w5100;
assign w6696 = ~w6694 & ~w6695;
assign w6697 = pi1454 & ~w5100;
assign w6698 = pi2177 & w5100;
assign w6699 = ~w6697 & ~w6698;
assign w6700 = pi1455 & ~w5100;
assign w6701 = pi2173 & w5100;
assign w6702 = ~w6700 & ~w6701;
assign w6703 = pi1456 & ~w5100;
assign w6704 = pi2194 & w5100;
assign w6705 = ~w6703 & ~w6704;
assign w6706 = pi1457 & ~w5100;
assign w6707 = pi2188 & w5100;
assign w6708 = ~w6706 & ~w6707;
assign w6709 = pi1458 & ~w5100;
assign w6710 = pi2184 & w5100;
assign w6711 = ~w6709 & ~w6710;
assign w6712 = pi1459 & ~w5100;
assign w6713 = pi2166 & w5100;
assign w6714 = ~w6712 & ~w6713;
assign w6715 = pi1460 & ~w5100;
assign w6716 = pi2192 & w5100;
assign w6717 = ~w6715 & ~w6716;
assign w6718 = ~pi0943 & w5104;
assign w6719 = pi1461 & ~w6718;
assign w6720 = pi2186 & w6718;
assign w6721 = ~w6719 & ~w6720;
assign w6722 = pi1462 & ~w6718;
assign w6723 = pi2183 & w6718;
assign w6724 = ~w6722 & ~w6723;
assign w6725 = pi1463 & ~w6718;
assign w6726 = pi2168 & w6718;
assign w6727 = ~w6725 & ~w6726;
assign w6728 = pi1464 & ~w6718;
assign w6729 = pi2174 & w6718;
assign w6730 = ~w6728 & ~w6729;
assign w6731 = pi1465 & ~w6718;
assign w6732 = pi2197 & w6718;
assign w6733 = ~w6731 & ~w6732;
assign w6734 = pi1466 & ~w6718;
assign w6735 = pi2196 & w6718;
assign w6736 = ~w6734 & ~w6735;
assign w6737 = pi1467 & ~w6718;
assign w6738 = pi2193 & w6718;
assign w6739 = ~w6737 & ~w6738;
assign w6740 = pi1468 & ~w6718;
assign w6741 = pi2189 & w6718;
assign w6742 = ~w6740 & ~w6741;
assign w6743 = pi1469 & ~w6718;
assign w6744 = pi2179 & w6718;
assign w6745 = ~w6743 & ~w6744;
assign w6746 = pi1470 & ~w6718;
assign w6747 = pi2198 & w6718;
assign w6748 = ~w6746 & ~w6747;
assign w6749 = pi1471 & ~w6718;
assign w6750 = pi2185 & w6718;
assign w6751 = ~w6749 & ~w6750;
assign w6752 = pi1472 & ~w6718;
assign w6753 = pi2187 & w6718;
assign w6754 = ~w6752 & ~w6753;
assign w6755 = pi1473 & ~w6718;
assign w6756 = pi2171 & w6718;
assign w6757 = ~w6755 & ~w6756;
assign w6758 = pi1474 & ~w6718;
assign w6759 = pi2169 & w6718;
assign w6760 = ~w6758 & ~w6759;
assign w6761 = pi1475 & ~w6718;
assign w6762 = pi2190 & w6718;
assign w6763 = ~w6761 & ~w6762;
assign w6764 = pi1476 & ~w6718;
assign w6765 = pi2181 & w6718;
assign w6766 = ~w6764 & ~w6765;
assign w6767 = pi1477 & ~w6718;
assign w6768 = pi2182 & w6718;
assign w6769 = ~w6767 & ~w6768;
assign w6770 = pi1478 & ~w6718;
assign w6771 = pi2175 & w6718;
assign w6772 = ~w6770 & ~w6771;
assign w6773 = pi1479 & ~w6718;
assign w6774 = pi2177 & w6718;
assign w6775 = ~w6773 & ~w6774;
assign w6776 = pi1480 & ~w6718;
assign w6777 = pi2173 & w6718;
assign w6778 = ~w6776 & ~w6777;
assign w6779 = pi1481 & ~w6718;
assign w6780 = pi2194 & w6718;
assign w6781 = ~w6779 & ~w6780;
assign w6782 = pi1482 & ~w6718;
assign w6783 = pi2188 & w6718;
assign w6784 = ~w6782 & ~w6783;
assign w6785 = pi1483 & ~w6718;
assign w6786 = pi2184 & w6718;
assign w6787 = ~w6785 & ~w6786;
assign w6788 = pi1484 & ~w6718;
assign w6789 = pi2166 & w6718;
assign w6790 = ~w6788 & ~w6789;
assign w6791 = pi1485 & ~w6718;
assign w6792 = pi2192 & w6718;
assign w6793 = ~w6791 & ~w6792;
assign w6794 = pi0943 & w5074;
assign w6795 = pi1486 & ~w6794;
assign w6796 = pi2186 & w6794;
assign w6797 = ~w6795 & ~w6796;
assign w6798 = pi1487 & ~w6794;
assign w6799 = pi2183 & w6794;
assign w6800 = ~w6798 & ~w6799;
assign w6801 = pi1488 & ~w6794;
assign w6802 = pi2168 & w6794;
assign w6803 = ~w6801 & ~w6802;
assign w6804 = pi1489 & ~w6794;
assign w6805 = pi2174 & w6794;
assign w6806 = ~w6804 & ~w6805;
assign w6807 = pi1490 & ~w6794;
assign w6808 = pi2197 & w6794;
assign w6809 = ~w6807 & ~w6808;
assign w6810 = pi1491 & ~w6794;
assign w6811 = pi2196 & w6794;
assign w6812 = ~w6810 & ~w6811;
assign w6813 = pi1492 & ~w6794;
assign w6814 = pi2193 & w6794;
assign w6815 = ~w6813 & ~w6814;
assign w6816 = pi1493 & ~w6794;
assign w6817 = pi2189 & w6794;
assign w6818 = ~w6816 & ~w6817;
assign w6819 = pi1494 & ~w6794;
assign w6820 = pi2198 & w6794;
assign w6821 = ~w6819 & ~w6820;
assign w6822 = pi1495 & ~w6794;
assign w6823 = pi2185 & w6794;
assign w6824 = ~w6822 & ~w6823;
assign w6825 = pi1496 & ~w6794;
assign w6826 = pi2187 & w6794;
assign w6827 = ~w6825 & ~w6826;
assign w6828 = pi1497 & ~w6794;
assign w6829 = pi2171 & w6794;
assign w6830 = ~w6828 & ~w6829;
assign w6831 = pi1498 & ~w6794;
assign w6832 = pi2169 & w6794;
assign w6833 = ~w6831 & ~w6832;
assign w6834 = pi1499 & ~w6794;
assign w6835 = pi2190 & w6794;
assign w6836 = ~w6834 & ~w6835;
assign w6837 = pi1500 & ~w6794;
assign w6838 = pi2181 & w6794;
assign w6839 = ~w6837 & ~w6838;
assign w6840 = pi1501 & ~w6794;
assign w6841 = pi2182 & w6794;
assign w6842 = ~w6840 & ~w6841;
assign w6843 = pi1502 & ~w6794;
assign w6844 = pi2175 & w6794;
assign w6845 = ~w6843 & ~w6844;
assign w6846 = pi1503 & ~w6794;
assign w6847 = pi2177 & w6794;
assign w6848 = ~w6846 & ~w6847;
assign w6849 = pi1504 & ~w6794;
assign w6850 = pi2173 & w6794;
assign w6851 = ~w6849 & ~w6850;
assign w6852 = pi1505 & ~w6794;
assign w6853 = pi2194 & w6794;
assign w6854 = ~w6852 & ~w6853;
assign w6855 = pi1506 & ~w6794;
assign w6856 = pi2188 & w6794;
assign w6857 = ~w6855 & ~w6856;
assign w6858 = pi1507 & ~w6794;
assign w6859 = pi2184 & w6794;
assign w6860 = ~w6858 & ~w6859;
assign w6861 = pi1508 & ~w6794;
assign w6862 = pi2166 & w6794;
assign w6863 = ~w6861 & ~w6862;
assign w6864 = pi1509 & ~w6794;
assign w6865 = pi2192 & w6794;
assign w6866 = ~w6864 & ~w6865;
assign w6867 = pi1510 & ~w5105;
assign w6868 = pi2186 & w5105;
assign w6869 = ~w6867 & ~w6868;
assign w6870 = pi1511 & ~w5105;
assign w6871 = pi2183 & w5105;
assign w6872 = ~w6870 & ~w6871;
assign w6873 = pi1512 & ~w5105;
assign w6874 = pi2168 & w5105;
assign w6875 = ~w6873 & ~w6874;
assign w6876 = pi1513 & ~w5105;
assign w6877 = pi2174 & w5105;
assign w6878 = ~w6876 & ~w6877;
assign w6879 = pi1514 & ~w5105;
assign w6880 = pi2197 & w5105;
assign w6881 = ~w6879 & ~w6880;
assign w6882 = pi1515 & ~w5105;
assign w6883 = pi2196 & w5105;
assign w6884 = ~w6882 & ~w6883;
assign w6885 = pi1516 & ~w5105;
assign w6886 = pi2193 & w5105;
assign w6887 = ~w6885 & ~w6886;
assign w6888 = pi1517 & ~w5105;
assign w6889 = pi2189 & w5105;
assign w6890 = ~w6888 & ~w6889;
assign w6891 = pi1518 & ~w5105;
assign w6892 = pi2198 & w5105;
assign w6893 = ~w6891 & ~w6892;
assign w6894 = pi1519 & ~w5105;
assign w6895 = pi2185 & w5105;
assign w6896 = ~w6894 & ~w6895;
assign w6897 = pi1520 & ~w5105;
assign w6898 = pi2187 & w5105;
assign w6899 = ~w6897 & ~w6898;
assign w6900 = pi1521 & ~w5105;
assign w6901 = pi2171 & w5105;
assign w6902 = ~w6900 & ~w6901;
assign w6903 = pi1522 & ~w5105;
assign w6904 = pi2169 & w5105;
assign w6905 = ~w6903 & ~w6904;
assign w6906 = pi1523 & ~w5105;
assign w6907 = pi2190 & w5105;
assign w6908 = ~w6906 & ~w6907;
assign w6909 = pi1524 & ~w5105;
assign w6910 = pi2181 & w5105;
assign w6911 = ~w6909 & ~w6910;
assign w6912 = pi1525 & ~w5105;
assign w6913 = pi2182 & w5105;
assign w6914 = ~w6912 & ~w6913;
assign w6915 = pi1526 & ~w5105;
assign w6916 = pi2175 & w5105;
assign w6917 = ~w6915 & ~w6916;
assign w6918 = pi1527 & ~w5105;
assign w6919 = pi2177 & w5105;
assign w6920 = ~w6918 & ~w6919;
assign w6921 = pi1528 & ~w5105;
assign w6922 = pi2173 & w5105;
assign w6923 = ~w6921 & ~w6922;
assign w6924 = pi1529 & ~w5105;
assign w6925 = pi2194 & w5105;
assign w6926 = ~w6924 & ~w6925;
assign w6927 = pi1530 & ~w5105;
assign w6928 = pi2188 & w5105;
assign w6929 = ~w6927 & ~w6928;
assign w6930 = pi1531 & ~w5105;
assign w6931 = pi2184 & w5105;
assign w6932 = ~w6930 & ~w6931;
assign w6933 = pi1532 & ~w5105;
assign w6934 = pi2166 & w5105;
assign w6935 = ~w6933 & ~w6934;
assign w6936 = pi1533 & ~w5105;
assign w6937 = pi2192 & w5105;
assign w6938 = ~w6936 & ~w6937;
assign w6939 = pi1534 & ~w5123;
assign w6940 = pi2195 & w5123;
assign w6941 = ~w6939 & ~w6940;
assign w6942 = pi1535 & ~w5166;
assign w6943 = pi2186 & w5166;
assign w6944 = ~w6942 & ~w6943;
assign w6945 = pi1536 & ~w5166;
assign w6946 = pi2172 & w5166;
assign w6947 = ~w6945 & ~w6946;
assign w6948 = pi1537 & ~w5166;
assign w6949 = pi2168 & w5166;
assign w6950 = ~w6948 & ~w6949;
assign w6951 = pi1538 & ~w5166;
assign w6952 = pi2174 & w5166;
assign w6953 = ~w6951 & ~w6952;
assign w6954 = pi1539 & ~w5166;
assign w6955 = pi2178 & w5166;
assign w6956 = ~w6954 & ~w6955;
assign w6957 = pi1540 & ~w5166;
assign w6958 = pi2196 & w5166;
assign w6959 = ~w6957 & ~w6958;
assign w6960 = pi1541 & ~w5166;
assign w6961 = pi2193 & w5166;
assign w6962 = ~w6960 & ~w6961;
assign w6963 = pi1542 & ~w5166;
assign w6964 = pi2189 & w5166;
assign w6965 = ~w6963 & ~w6964;
assign w6966 = pi1543 & ~w5166;
assign w6967 = pi2179 & w5166;
assign w6968 = ~w6966 & ~w6967;
assign w6969 = pi1544 & ~w5166;
assign w6970 = pi2198 & w5166;
assign w6971 = ~w6969 & ~w6970;
assign w6972 = pi1545 & ~w5166;
assign w6973 = pi2185 & w5166;
assign w6974 = ~w6972 & ~w6973;
assign w6975 = pi1546 & ~w5166;
assign w6976 = pi2176 & w5166;
assign w6977 = ~w6975 & ~w6976;
assign w6978 = pi1547 & ~w5166;
assign w6979 = pi2171 & w5166;
assign w6980 = ~w6978 & ~w6979;
assign w6981 = pi1548 & ~w5166;
assign w6982 = pi2169 & w5166;
assign w6983 = ~w6981 & ~w6982;
assign w6984 = pi1549 & ~w5166;
assign w6985 = pi2170 & w5166;
assign w6986 = ~w6984 & ~w6985;
assign w6987 = pi1550 & ~w5166;
assign w6988 = pi2181 & w5166;
assign w6989 = ~w6987 & ~w6988;
assign w6990 = pi1551 & ~w5166;
assign w6991 = pi2182 & w5166;
assign w6992 = ~w6990 & ~w6991;
assign w6993 = pi1552 & ~w5166;
assign w6994 = pi2191 & w5166;
assign w6995 = ~w6993 & ~w6994;
assign w6996 = pi1553 & ~w5166;
assign w6997 = pi2177 & w5166;
assign w6998 = ~w6996 & ~w6997;
assign w6999 = pi1554 & ~w5166;
assign w7000 = pi2173 & w5166;
assign w7001 = ~w6999 & ~w7000;
assign w7002 = pi1555 & ~w5166;
assign w7003 = pi2167 & w5166;
assign w7004 = ~w7002 & ~w7003;
assign w7005 = pi1556 & ~w5166;
assign w7006 = pi2188 & w5166;
assign w7007 = ~w7005 & ~w7006;
assign w7008 = pi1557 & ~w5166;
assign w7009 = pi2184 & w5166;
assign w7010 = ~w7008 & ~w7009;
assign w7011 = pi1558 & ~w5166;
assign w7012 = pi2195 & w5166;
assign w7013 = ~w7011 & ~w7012;
assign w7014 = pi1559 & ~w5166;
assign w7015 = pi2192 & w5166;
assign w7016 = ~w7014 & ~w7015;
assign w7017 = pi1560 & ~w5647;
assign w7018 = pi2186 & w5647;
assign w7019 = ~w7017 & ~w7018;
assign w7020 = pi1561 & ~w5647;
assign w7021 = pi2172 & w5647;
assign w7022 = ~w7020 & ~w7021;
assign w7023 = pi1562 & ~w5647;
assign w7024 = pi2168 & w5647;
assign w7025 = ~w7023 & ~w7024;
assign w7026 = pi1563 & ~w5647;
assign w7027 = pi2174 & w5647;
assign w7028 = ~w7026 & ~w7027;
assign w7029 = pi1564 & ~w5647;
assign w7030 = pi2178 & w5647;
assign w7031 = ~w7029 & ~w7030;
assign w7032 = pi1565 & ~w5647;
assign w7033 = pi2196 & w5647;
assign w7034 = ~w7032 & ~w7033;
assign w7035 = pi1566 & ~w5647;
assign w7036 = pi2193 & w5647;
assign w7037 = ~w7035 & ~w7036;
assign w7038 = pi1567 & ~w5647;
assign w7039 = pi2179 & w5647;
assign w7040 = ~w7038 & ~w7039;
assign w7041 = pi1568 & ~w5647;
assign w7042 = pi2198 & w5647;
assign w7043 = ~w7041 & ~w7042;
assign w7044 = pi1569 & ~w5647;
assign w7045 = pi2185 & w5647;
assign w7046 = ~w7044 & ~w7045;
assign w7047 = pi1570 & ~w5647;
assign w7048 = pi2176 & w5647;
assign w7049 = ~w7047 & ~w7048;
assign w7050 = pi1571 & ~w5647;
assign w7051 = pi2171 & w5647;
assign w7052 = ~w7050 & ~w7051;
assign w7053 = pi1572 & ~w5647;
assign w7054 = pi2169 & w5647;
assign w7055 = ~w7053 & ~w7054;
assign w7056 = pi1573 & ~w5647;
assign w7057 = pi2170 & w5647;
assign w7058 = ~w7056 & ~w7057;
assign w7059 = pi1574 & ~w5647;
assign w7060 = pi2181 & w5647;
assign w7061 = ~w7059 & ~w7060;
assign w7062 = pi1575 & ~w5647;
assign w7063 = pi2182 & w5647;
assign w7064 = ~w7062 & ~w7063;
assign w7065 = pi1576 & ~w5647;
assign w7066 = pi2191 & w5647;
assign w7067 = ~w7065 & ~w7066;
assign w7068 = pi1577 & ~w5647;
assign w7069 = pi2177 & w5647;
assign w7070 = ~w7068 & ~w7069;
assign w7071 = pi1578 & ~w5647;
assign w7072 = pi2173 & w5647;
assign w7073 = ~w7071 & ~w7072;
assign w7074 = pi1579 & ~w5647;
assign w7075 = pi2167 & w5647;
assign w7076 = ~w7074 & ~w7075;
assign w7077 = pi1580 & ~w5647;
assign w7078 = pi2188 & w5647;
assign w7079 = ~w7077 & ~w7078;
assign w7080 = pi1581 & ~w5647;
assign w7081 = pi2184 & w5647;
assign w7082 = ~w7080 & ~w7081;
assign w7083 = pi1582 & ~w5647;
assign w7084 = pi2195 & w5647;
assign w7085 = ~w7083 & ~w7084;
assign w7086 = pi1583 & ~w5647;
assign w7087 = pi2192 & w5647;
assign w7088 = ~w7086 & ~w7087;
assign w7089 = pi1584 & ~w5132;
assign w7090 = pi2186 & w5132;
assign w7091 = ~w7089 & ~w7090;
assign w7092 = pi1585 & ~w5132;
assign w7093 = pi2172 & w5132;
assign w7094 = ~w7092 & ~w7093;
assign w7095 = pi1586 & ~w5132;
assign w7096 = pi2168 & w5132;
assign w7097 = ~w7095 & ~w7096;
assign w7098 = pi1587 & ~w5132;
assign w7099 = pi2174 & w5132;
assign w7100 = ~w7098 & ~w7099;
assign w7101 = pi1588 & ~w5132;
assign w7102 = pi2178 & w5132;
assign w7103 = ~w7101 & ~w7102;
assign w7104 = pi1589 & ~w5132;
assign w7105 = pi2196 & w5132;
assign w7106 = ~w7104 & ~w7105;
assign w7107 = pi1590 & ~w5132;
assign w7108 = pi2193 & w5132;
assign w7109 = ~w7107 & ~w7108;
assign w7110 = pi1591 & ~w5132;
assign w7111 = pi2179 & w5132;
assign w7112 = ~w7110 & ~w7111;
assign w7113 = pi1592 & ~w5132;
assign w7114 = pi2198 & w5132;
assign w7115 = ~w7113 & ~w7114;
assign w7116 = pi1593 & ~w5132;
assign w7117 = pi2185 & w5132;
assign w7118 = ~w7116 & ~w7117;
assign w7119 = pi1594 & ~w5252;
assign w7120 = pi2185 & w5252;
assign w7121 = ~w7119 & ~w7120;
assign w7122 = pi1595 & ~w5132;
assign w7123 = pi2176 & w5132;
assign w7124 = ~w7122 & ~w7123;
assign w7125 = pi1596 & ~w5132;
assign w7126 = pi2171 & w5132;
assign w7127 = ~w7125 & ~w7126;
assign w7128 = pi1597 & ~w5132;
assign w7129 = pi2169 & w5132;
assign w7130 = ~w7128 & ~w7129;
assign w7131 = pi1598 & ~w5132;
assign w7132 = pi2170 & w5132;
assign w7133 = ~w7131 & ~w7132;
assign w7134 = pi1599 & ~w5132;
assign w7135 = pi2181 & w5132;
assign w7136 = ~w7134 & ~w7135;
assign w7137 = pi1600 & ~w5132;
assign w7138 = pi2182 & w5132;
assign w7139 = ~w7137 & ~w7138;
assign w7140 = pi1601 & ~w5132;
assign w7141 = pi2191 & w5132;
assign w7142 = ~w7140 & ~w7141;
assign w7143 = pi1602 & ~w5132;
assign w7144 = pi2177 & w5132;
assign w7145 = ~w7143 & ~w7144;
assign w7146 = pi1603 & ~w5132;
assign w7147 = pi2173 & w5132;
assign w7148 = ~w7146 & ~w7147;
assign w7149 = pi1604 & ~w5132;
assign w7150 = pi2167 & w5132;
assign w7151 = ~w7149 & ~w7150;
assign w7152 = pi1605 & ~w5132;
assign w7153 = pi2188 & w5132;
assign w7154 = ~w7152 & ~w7153;
assign w7155 = pi1606 & ~w5132;
assign w7156 = pi2184 & w5132;
assign w7157 = ~w7155 & ~w7156;
assign w7158 = pi1607 & ~w5132;
assign w7159 = pi2195 & w5132;
assign w7160 = ~w7158 & ~w7159;
assign w7161 = pi1608 & ~w5132;
assign w7162 = pi2192 & w5132;
assign w7163 = ~w7161 & ~w7162;
assign w7164 = pi1609 & ~w5152;
assign w7165 = pi2186 & w5152;
assign w7166 = ~w7164 & ~w7165;
assign w7167 = pi1610 & ~w5152;
assign w7168 = pi2172 & w5152;
assign w7169 = ~w7167 & ~w7168;
assign w7170 = pi1611 & ~w5152;
assign w7171 = pi2168 & w5152;
assign w7172 = ~w7170 & ~w7171;
assign w7173 = pi1612 & ~w5152;
assign w7174 = pi2174 & w5152;
assign w7175 = ~w7173 & ~w7174;
assign w7176 = pi1613 & ~w5152;
assign w7177 = pi2178 & w5152;
assign w7178 = ~w7176 & ~w7177;
assign w7179 = pi1614 & ~w5152;
assign w7180 = pi2196 & w5152;
assign w7181 = ~w7179 & ~w7180;
assign w7182 = pi1615 & ~w5152;
assign w7183 = pi2193 & w5152;
assign w7184 = ~w7182 & ~w7183;
assign w7185 = pi1616 & ~w5152;
assign w7186 = pi2179 & w5152;
assign w7187 = ~w7185 & ~w7186;
assign w7188 = pi1617 & ~w5152;
assign w7189 = pi2198 & w5152;
assign w7190 = ~w7188 & ~w7189;
assign w7191 = pi1618 & ~w5152;
assign w7192 = pi2185 & w5152;
assign w7193 = ~w7191 & ~w7192;
assign w7194 = pi1619 & ~w5152;
assign w7195 = pi2176 & w5152;
assign w7196 = ~w7194 & ~w7195;
assign w7197 = pi1620 & ~w5152;
assign w7198 = pi2171 & w5152;
assign w7199 = ~w7197 & ~w7198;
assign w7200 = pi1621 & ~w5152;
assign w7201 = pi2169 & w5152;
assign w7202 = ~w7200 & ~w7201;
assign w7203 = pi1622 & ~w5152;
assign w7204 = pi2170 & w5152;
assign w7205 = ~w7203 & ~w7204;
assign w7206 = pi1623 & ~w5422;
assign w7207 = pi2186 & w5422;
assign w7208 = ~w7206 & ~w7207;
assign w7209 = pi1624 & ~w5152;
assign w7210 = pi2181 & w5152;
assign w7211 = ~w7209 & ~w7210;
assign w7212 = pi1625 & ~w5422;
assign w7213 = pi2183 & w5422;
assign w7214 = ~w7212 & ~w7213;
assign w7215 = pi1626 & ~w5152;
assign w7216 = pi2175 & w5152;
assign w7217 = ~w7215 & ~w7216;
assign w7218 = pi1627 & ~w5152;
assign w7219 = pi2191 & w5152;
assign w7220 = ~w7218 & ~w7219;
assign w7221 = pi1628 & ~w5152;
assign w7222 = pi2177 & w5152;
assign w7223 = ~w7221 & ~w7222;
assign w7224 = pi1629 & ~w5152;
assign w7225 = pi2173 & w5152;
assign w7226 = ~w7224 & ~w7225;
assign w7227 = pi1630 & ~w5422;
assign w7228 = pi2168 & w5422;
assign w7229 = ~w7227 & ~w7228;
assign w7230 = pi1631 & ~w5152;
assign w7231 = pi2167 & w5152;
assign w7232 = ~w7230 & ~w7231;
assign w7233 = pi1632 & ~w5422;
assign w7234 = pi2174 & w5422;
assign w7235 = ~w7233 & ~w7234;
assign w7236 = pi1633 & ~w5152;
assign w7237 = pi2188 & w5152;
assign w7238 = ~w7236 & ~w7237;
assign w7239 = pi1634 & ~w5422;
assign w7240 = pi2197 & w5422;
assign w7241 = ~w7239 & ~w7240;
assign w7242 = pi1635 & ~w5152;
assign w7243 = pi2166 & w5152;
assign w7244 = ~w7242 & ~w7243;
assign w7245 = pi1636 & ~w5152;
assign w7246 = pi2195 & w5152;
assign w7247 = ~w7245 & ~w7246;
assign w7248 = pi1637 & ~w5152;
assign w7249 = pi2192 & w5152;
assign w7250 = ~w7248 & ~w7249;
assign w7251 = pi1638 & ~w5385;
assign w7252 = pi2186 & w5385;
assign w7253 = ~w7251 & ~w7252;
assign w7254 = pi1639 & ~w5422;
assign w7255 = pi2196 & w5422;
assign w7256 = ~w7254 & ~w7255;
assign w7257 = pi1640 & ~w5385;
assign w7258 = pi2183 & w5385;
assign w7259 = ~w7257 & ~w7258;
assign w7260 = pi1641 & ~w5385;
assign w7261 = pi2172 & w5385;
assign w7262 = ~w7260 & ~w7261;
assign w7263 = pi1642 & ~w5422;
assign w7264 = pi2193 & w5422;
assign w7265 = ~w7263 & ~w7264;
assign w7266 = pi1643 & ~w5385;
assign w7267 = pi2168 & w5385;
assign w7268 = ~w7266 & ~w7267;
assign w7269 = pi1644 & ~w5422;
assign w7270 = pi2189 & w5422;
assign w7271 = ~w7269 & ~w7270;
assign w7272 = pi1645 & ~w5385;
assign w7273 = pi2197 & w5385;
assign w7274 = ~w7272 & ~w7273;
assign w7275 = pi1646 & ~w5385;
assign w7276 = pi2178 & w5385;
assign w7277 = ~w7275 & ~w7276;
assign w7278 = pi1647 & ~w5385;
assign w7279 = pi2196 & w5385;
assign w7280 = ~w7278 & ~w7279;
assign w7281 = pi1648 & ~w5385;
assign w7282 = pi2193 & w5385;
assign w7283 = ~w7281 & ~w7282;
assign w7284 = pi1649 & ~w5422;
assign w7285 = pi2198 & w5422;
assign w7286 = ~w7284 & ~w7285;
assign w7287 = pi1650 & ~w5385;
assign w7288 = pi2179 & w5385;
assign w7289 = ~w7287 & ~w7288;
assign w7290 = pi1651 & ~w5422;
assign w7291 = pi2185 & w5422;
assign w7292 = ~w7290 & ~w7291;
assign w7293 = pi1652 & ~w5385;
assign w7294 = pi2198 & w5385;
assign w7295 = ~w7293 & ~w7294;
assign w7296 = pi1653 & ~w5422;
assign w7297 = pi2187 & w5422;
assign w7298 = ~w7296 & ~w7297;
assign w7299 = pi1654 & ~w5385;
assign w7300 = pi2187 & w5385;
assign w7301 = ~w7299 & ~w7300;
assign w7302 = pi1655 & ~w5385;
assign w7303 = pi2176 & w5385;
assign w7304 = ~w7302 & ~w7303;
assign w7305 = pi1656 & ~w5385;
assign w7306 = pi2171 & w5385;
assign w7307 = ~w7305 & ~w7306;
assign w7308 = pi1657 & ~w5385;
assign w7309 = pi2169 & w5385;
assign w7310 = ~w7308 & ~w7309;
assign w7311 = pi1658 & ~w5422;
assign w7312 = pi2171 & w5422;
assign w7313 = ~w7311 & ~w7312;
assign w7314 = pi1659 & ~w5385;
assign w7315 = pi2170 & w5385;
assign w7316 = ~w7314 & ~w7315;
assign w7317 = pi1660 & ~w5422;
assign w7318 = pi2169 & w5422;
assign w7319 = ~w7317 & ~w7318;
assign w7320 = pi1661 & ~w5385;
assign w7321 = pi2181 & w5385;
assign w7322 = ~w7320 & ~w7321;
assign w7323 = pi1662 & ~w5422;
assign w7324 = pi2190 & w5422;
assign w7325 = ~w7323 & ~w7324;
assign w7326 = pi1663 & ~w5385;
assign w7327 = pi2175 & w5385;
assign w7328 = ~w7326 & ~w7327;
assign w7329 = pi1664 & ~w5385;
assign w7330 = pi2191 & w5385;
assign w7331 = ~w7329 & ~w7330;
assign w7332 = pi1665 & ~w5385;
assign w7333 = pi2177 & w5385;
assign w7334 = ~w7332 & ~w7333;
assign w7335 = pi1666 & ~w5385;
assign w7336 = pi2173 & w5385;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = pi1667 & ~w5422;
assign w7339 = pi2181 & w5422;
assign w7340 = ~w7338 & ~w7339;
assign w7341 = pi1668 & ~w5190;
assign w7342 = pi2186 & w5190;
assign w7343 = ~w7341 & ~w7342;
assign w7344 = pi1669 & ~w5190;
assign w7345 = pi2183 & w5190;
assign w7346 = ~w7344 & ~w7345;
assign w7347 = pi1670 & ~w5190;
assign w7348 = pi2172 & w5190;
assign w7349 = ~w7347 & ~w7348;
assign w7350 = pi1671 & ~w5190;
assign w7351 = pi2178 & w5190;
assign w7352 = ~w7350 & ~w7351;
assign w7353 = pi1672 & ~w5190;
assign w7354 = pi2189 & w5190;
assign w7355 = ~w7353 & ~w7354;
assign w7356 = pi1673 & ~w5190;
assign w7357 = pi2198 & w5190;
assign w7358 = ~w7356 & ~w7357;
assign w7359 = pi1674 & ~w5190;
assign w7360 = pi2187 & w5190;
assign w7361 = ~w7359 & ~w7360;
assign w7362 = pi1675 & ~w5190;
assign w7363 = pi2190 & w5190;
assign w7364 = ~w7362 & ~w7363;
assign w7365 = pi1676 & ~w5190;
assign w7366 = pi2181 & w5190;
assign w7367 = ~w7365 & ~w7366;
assign w7368 = pi1677 & ~w5190;
assign w7369 = pi2182 & w5190;
assign w7370 = ~w7368 & ~w7369;
assign w7371 = pi1678 & ~w5190;
assign w7372 = pi2170 & w5190;
assign w7373 = ~w7371 & ~w7372;
assign w7374 = pi1679 & ~w5190;
assign w7375 = pi2191 & w5190;
assign w7376 = ~w7374 & ~w7375;
assign w7377 = pi1680 & ~w5190;
assign w7378 = pi2175 & w5190;
assign w7379 = ~w7377 & ~w7378;
assign w7380 = pi1681 & ~w5190;
assign w7381 = pi2194 & w5190;
assign w7382 = ~w7380 & ~w7381;
assign w7383 = pi1682 & ~w5190;
assign w7384 = pi2188 & w5190;
assign w7385 = ~w7383 & ~w7384;
assign w7386 = pi1683 & ~w5190;
assign w7387 = pi2195 & w5190;
assign w7388 = ~w7386 & ~w7387;
assign w7389 = pi1684 & ~w5221;
assign w7390 = pi2183 & w5221;
assign w7391 = ~w7389 & ~w7390;
assign w7392 = pi1685 & ~w5221;
assign w7393 = pi2172 & w5221;
assign w7394 = ~w7392 & ~w7393;
assign w7395 = pi1686 & ~w5221;
assign w7396 = pi2178 & w5221;
assign w7397 = ~w7395 & ~w7396;
assign w7398 = pi1687 & ~w5221;
assign w7399 = pi2189 & w5221;
assign w7400 = ~w7398 & ~w7399;
assign w7401 = pi1688 & ~w5221;
assign w7402 = pi2198 & w5221;
assign w7403 = ~w7401 & ~w7402;
assign w7404 = pi1689 & ~w5221;
assign w7405 = pi2187 & w5221;
assign w7406 = ~w7404 & ~w7405;
assign w7407 = pi1690 & ~w5729;
assign w7408 = pi2195 & w5729;
assign w7409 = ~w7407 & ~w7408;
assign w7410 = pi1691 & ~w5221;
assign w7411 = pi2170 & w5221;
assign w7412 = ~w7410 & ~w7411;
assign w7413 = pi1692 & ~w5221;
assign w7414 = pi2181 & w5221;
assign w7415 = ~w7413 & ~w7414;
assign w7416 = pi1693 & ~w5221;
assign w7417 = pi2190 & w5221;
assign w7418 = ~w7416 & ~w7417;
assign w7419 = pi1694 & ~w5221;
assign w7420 = pi2191 & w5221;
assign w7421 = ~w7419 & ~w7420;
assign w7422 = pi1695 & ~w5221;
assign w7423 = pi2175 & w5221;
assign w7424 = ~w7422 & ~w7423;
assign w7425 = pi1696 & ~w5221;
assign w7426 = pi2194 & w5221;
assign w7427 = ~w7425 & ~w7426;
assign w7428 = pi1697 & ~w5221;
assign w7429 = pi2188 & w5221;
assign w7430 = ~w7428 & ~w7429;
assign w7431 = pi1698 & ~w5221;
assign w7432 = pi2195 & w5221;
assign w7433 = ~w7431 & ~w7432;
assign w7434 = pi1699 & ~w5252;
assign w7435 = pi2183 & w5252;
assign w7436 = ~w7434 & ~w7435;
assign w7437 = pi1700 & ~w5252;
assign w7438 = pi2172 & w5252;
assign w7439 = ~w7437 & ~w7438;
assign w7440 = pi1701 & ~w5252;
assign w7441 = pi2178 & w5252;
assign w7442 = ~w7440 & ~w7441;
assign w7443 = pi1702 & ~w5166;
assign w7444 = pi2187 & w5166;
assign w7445 = ~w7443 & ~w7444;
assign w7446 = pi1703 & ~w5252;
assign w7447 = pi2189 & w5252;
assign w7448 = ~w7446 & ~w7447;
assign w7449 = pi1704 & ~w5252;
assign w7450 = pi2198 & w5252;
assign w7451 = ~w7449 & ~w7450;
assign w7452 = pi1705 & ~w5252;
assign w7453 = pi2187 & w5252;
assign w7454 = ~w7452 & ~w7453;
assign w7455 = pi1706 & ~w5252;
assign w7456 = pi2170 & w5252;
assign w7457 = ~w7455 & ~w7456;
assign w7458 = pi1707 & ~w5252;
assign w7459 = pi2181 & w5252;
assign w7460 = ~w7458 & ~w7459;
assign w7461 = pi1708 & ~w5252;
assign w7462 = pi2190 & w5252;
assign w7463 = ~w7461 & ~w7462;
assign w7464 = pi1709 & ~w5252;
assign w7465 = pi2191 & w5252;
assign w7466 = ~w7464 & ~w7465;
assign w7467 = pi1710 & ~w5252;
assign w7468 = pi2175 & w5252;
assign w7469 = ~w7467 & ~w7468;
assign w7470 = pi1711 & ~w5252;
assign w7471 = pi2194 & w5252;
assign w7472 = ~w7470 & ~w7471;
assign w7473 = pi1712 & ~w5252;
assign w7474 = pi2188 & w5252;
assign w7475 = ~w7473 & ~w7474;
assign w7476 = pi1713 & ~w5252;
assign w7477 = pi2195 & w5252;
assign w7478 = ~w7476 & ~w7477;
assign w7479 = pi1714 & ~w5284;
assign w7480 = pi2183 & w5284;
assign w7481 = ~w7479 & ~w7480;
assign w7482 = pi1715 & ~w5284;
assign w7483 = pi2172 & w5284;
assign w7484 = ~w7482 & ~w7483;
assign w7485 = pi1716 & ~w5284;
assign w7486 = pi2178 & w5284;
assign w7487 = ~w7485 & ~w7486;
assign w7488 = pi1717 & ~w5284;
assign w7489 = pi2189 & w5284;
assign w7490 = ~w7488 & ~w7489;
assign w7491 = pi1718 & ~w5284;
assign w7492 = pi2198 & w5284;
assign w7493 = ~w7491 & ~w7492;
assign w7494 = pi1719 & ~w5284;
assign w7495 = pi2187 & w5284;
assign w7496 = ~w7494 & ~w7495;
assign w7497 = pi1720 & ~w5284;
assign w7498 = pi2190 & w5284;
assign w7499 = ~w7497 & ~w7498;
assign w7500 = pi1721 & ~w5284;
assign w7501 = pi2181 & w5284;
assign w7502 = ~w7500 & ~w7501;
assign w7503 = pi1722 & ~w5284;
assign w7504 = pi2182 & w5284;
assign w7505 = ~w7503 & ~w7504;
assign w7506 = pi1723 & ~w5284;
assign w7507 = pi2170 & w5284;
assign w7508 = ~w7506 & ~w7507;
assign w7509 = pi1724 & ~w5284;
assign w7510 = pi2191 & w5284;
assign w7511 = ~w7509 & ~w7510;
assign w7512 = pi1725 & ~w5284;
assign w7513 = pi2175 & w5284;
assign w7514 = ~w7512 & ~w7513;
assign w7515 = pi1726 & ~w5284;
assign w7516 = pi2194 & w5284;
assign w7517 = ~w7515 & ~w7516;
assign w7518 = pi1727 & ~w5284;
assign w7519 = pi2188 & w5284;
assign w7520 = ~w7518 & ~w7519;
assign w7521 = pi1728 & ~w5284;
assign w7522 = pi2195 & w5284;
assign w7523 = ~w7521 & ~w7522;
assign w7524 = pi1729 & ~w5315;
assign w7525 = pi2183 & w5315;
assign w7526 = ~w7524 & ~w7525;
assign w7527 = pi1730 & ~w5326;
assign w7528 = pi2183 & w5326;
assign w7529 = ~w7527 & ~w7528;
assign w7530 = pi1731 & ~w5326;
assign w7531 = pi2174 & w5326;
assign w7532 = ~w7530 & ~w7531;
assign w7533 = pi1732 & ~w5315;
assign w7534 = pi2189 & w5315;
assign w7535 = ~w7533 & ~w7534;
assign w7536 = pi1733 & ~w5326;
assign w7537 = pi2197 & w5326;
assign w7538 = ~w7536 & ~w7537;
assign w7539 = pi1734 & ~w5315;
assign w7540 = pi2179 & w5315;
assign w7541 = ~w7539 & ~w7540;
assign w7542 = pi1735 & ~w5326;
assign w7543 = pi2189 & w5326;
assign w7544 = ~w7542 & ~w7543;
assign w7545 = pi1736 & ~w5326;
assign w7546 = pi2179 & w5326;
assign w7547 = ~w7545 & ~w7546;
assign w7548 = pi1737 & ~w5315;
assign w7549 = pi2185 & w5315;
assign w7550 = ~w7548 & ~w7549;
assign w7551 = pi1738 & ~w5326;
assign w7552 = pi2185 & w5326;
assign w7553 = ~w7551 & ~w7552;
assign w7554 = pi1739 & ~w5326;
assign w7555 = pi2187 & w5326;
assign w7556 = ~w7554 & ~w7555;
assign w7557 = pi1740 & ~w5315;
assign w7558 = pi2176 & w5315;
assign w7559 = ~w7557 & ~w7558;
assign w7560 = pi1741 & ~w5326;
assign w7561 = pi2171 & w5326;
assign w7562 = ~w7560 & ~w7561;
assign w7563 = pi1742 & ~w5326;
assign w7564 = pi2169 & w5326;
assign w7565 = ~w7563 & ~w7564;
assign w7566 = pi1743 & ~w5326;
assign w7567 = pi2190 & w5326;
assign w7568 = ~w7566 & ~w7567;
assign w7569 = pi1744 & ~w5315;
assign w7570 = pi2169 & w5315;
assign w7571 = ~w7569 & ~w7570;
assign w7572 = pi1745 & ~w5315;
assign w7573 = pi2190 & w5315;
assign w7574 = ~w7572 & ~w7573;
assign w7575 = pi1746 & ~w5315;
assign w7576 = pi2170 & w5315;
assign w7577 = ~w7575 & ~w7576;
assign w7578 = pi1747 & ~w5315;
assign w7579 = pi2182 & w5315;
assign w7580 = ~w7578 & ~w7579;
assign w7581 = pi1748 & ~w5326;
assign w7582 = pi2166 & w5326;
assign w7583 = ~w7581 & ~w7582;
assign w7584 = pi1749 & ~w5326;
assign w7585 = pi2195 & w5326;
assign w7586 = ~w7584 & ~w7585;
assign w7587 = pi1750 & ~w5326;
assign w7588 = pi2184 & w5326;
assign w7589 = ~w7587 & ~w7588;
assign w7590 = pi1751 & ~w5326;
assign w7591 = pi2192 & w5326;
assign w7592 = ~w7590 & ~w7591;
assign w7593 = pi1752 & ~w5315;
assign w7594 = pi2177 & w5315;
assign w7595 = ~w7593 & ~w7594;
assign w7596 = pi1753 & ~w5315;
assign w7597 = pi2194 & w5315;
assign w7598 = ~w7596 & ~w7597;
assign w7599 = pi1754 & ~w5315;
assign w7600 = pi2195 & w5315;
assign w7601 = ~w7599 & ~w7600;
assign w7602 = pi1755 & ~w5166;
assign w7603 = pi2183 & w5166;
assign w7604 = ~w7602 & ~w7603;
assign w7605 = pi1756 & ~w5378;
assign w7606 = ~pi2166 & w5378;
assign w7607 = ~w7605 & ~w7606;
assign w7608 = pi1757 & ~w6794;
assign w7609 = pi2176 & w6794;
assign w7610 = ~w7608 & ~w7609;
assign w7611 = pi1758 & ~w5252;
assign w7612 = pi2186 & w5252;
assign w7613 = ~w7611 & ~w7612;
assign w7614 = pi1759 & ~w5105;
assign w7615 = pi2167 & w5105;
assign w7616 = ~w7614 & ~w7615;
assign w7617 = pi1760 & ~w5729;
assign w7618 = pi2170 & w5729;
assign w7619 = ~w7617 & ~w7618;
assign w7620 = pi1761 & ~w5105;
assign w7621 = pi2191 & w5105;
assign w7622 = ~w7620 & ~w7621;
assign w7623 = pi1762 & ~w5406;
assign w7624 = pi2176 & w5406;
assign w7625 = ~w7623 & ~w7624;
assign w7626 = pi1763 & ~w5105;
assign w7627 = pi2170 & w5105;
assign w7628 = ~w7626 & ~w7627;
assign w7629 = pi1764 & ~w5105;
assign w7630 = pi2176 & w5105;
assign w7631 = ~w7629 & ~w7630;
assign w7632 = pi1765 & ~w5105;
assign w7633 = pi2178 & w5105;
assign w7634 = ~w7632 & ~w7633;
assign w7635 = pi1766 & ~w5221;
assign w7636 = pi2184 & w5221;
assign w7637 = ~w7635 & ~w7636;
assign w7638 = pi1767 & ~w5105;
assign w7639 = pi2179 & w5105;
assign w7640 = ~w7638 & ~w7639;
assign w7641 = pi1769 & ~w5221;
assign w7642 = pi2177 & w5221;
assign w7643 = ~w7641 & ~w7642;
assign w7644 = pi1770 & ~w5221;
assign w7645 = pi2171 & w5221;
assign w7646 = ~w7644 & ~w7645;
assign w7647 = pi1771 & ~w5378;
assign w7648 = pi2189 & w5378;
assign w7649 = ~w7647 & ~w7648;
assign w7650 = pi1772 & ~w6794;
assign w7651 = pi2167 & w6794;
assign w7652 = ~w7650 & ~w7651;
assign w7653 = pi1773 & ~w5105;
assign w7654 = pi2172 & w5105;
assign w7655 = ~w7653 & ~w7654;
assign w7656 = pi1774 & ~w6794;
assign w7657 = pi2195 & w6794;
assign w7658 = ~w7656 & ~w7657;
assign w7659 = pi1775 & ~w6794;
assign w7660 = pi2191 & w6794;
assign w7661 = ~w7659 & ~w7660;
assign w7662 = pi1776 & ~w5315;
assign w7663 = pi2192 & w5315;
assign w7664 = ~w7662 & ~w7663;
assign w7665 = pi1777 & ~w5406;
assign w7666 = pi2170 & w5406;
assign w7667 = ~w7665 & ~w7666;
assign w7668 = pi1778 & ~w5221;
assign w7669 = pi2182 & w5221;
assign w7670 = ~w7668 & ~w7669;
assign w7671 = pi1779 & ~w5729;
assign w7672 = pi2194 & w5729;
assign w7673 = ~w7671 & ~w7672;
assign w7674 = pi1780 & ~w6794;
assign w7675 = pi2170 & w6794;
assign w7676 = ~w7674 & ~w7675;
assign w7677 = pi1781 & ~w5315;
assign w7678 = pi2167 & w5315;
assign w7679 = ~w7677 & ~w7678;
assign w7680 = pi1782 & ~w5221;
assign w7681 = pi2185 & w5221;
assign w7682 = ~w7680 & ~w7681;
assign w7683 = pi1783 & ~w5326;
assign w7684 = pi2173 & w5326;
assign w7685 = ~w7683 & ~w7684;
assign w7686 = pi1784 & ~w6794;
assign w7687 = pi2178 & w6794;
assign w7688 = ~w7686 & ~w7687;
assign w7689 = pi1785 & ~w6718;
assign w7690 = pi2178 & w6718;
assign w7691 = ~w7689 & ~w7690;
assign w7692 = pi1786 & ~w6794;
assign w7693 = pi2179 & w6794;
assign w7694 = ~w7692 & ~w7693;
assign w7695 = pi1787 & ~w6794;
assign w7696 = pi2172 & w6794;
assign w7697 = ~w7695 & ~w7696;
assign w7698 = pi1788 & ~w5221;
assign w7699 = pi2193 & w5221;
assign w7700 = ~w7698 & ~w7699;
assign w7701 = pi1789 & ~w5406;
assign w7702 = pi2179 & w5406;
assign w7703 = ~w7701 & ~w7702;
assign w7704 = pi1790 & ~w5221;
assign w7705 = pi2168 & w5221;
assign w7706 = ~w7704 & ~w7705;
assign w7707 = pi1791 & ~w6718;
assign w7708 = pi2170 & w6718;
assign w7709 = ~w7707 & ~w7708;
assign w7710 = pi1792 & ~w5190;
assign w7711 = pi2184 & w5190;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = pi1793 & ~w6718;
assign w7714 = pi2167 & w6718;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = pi1794 & ~w6718;
assign w7717 = pi2195 & w6718;
assign w7718 = ~w7716 & ~w7717;
assign w7719 = pi1795 & ~w6718;
assign w7720 = pi2191 & w6718;
assign w7721 = ~w7719 & ~w7720;
assign w7722 = pi1796 & ~w5221;
assign w7723 = pi2186 & w5221;
assign w7724 = ~w7722 & ~w7723;
assign w7725 = pi1797 & ~w6718;
assign w7726 = pi2176 & w6718;
assign w7727 = ~w7725 & ~w7726;
assign w7728 = pi1798 & ~w5326;
assign w7729 = pi2194 & w5326;
assign w7730 = ~w7728 & ~w7729;
assign w7731 = pi1799 & ~w5190;
assign w7732 = pi2177 & w5190;
assign w7733 = ~w7731 & ~w7732;
assign w7734 = pi1800 & ~w5326;
assign w7735 = pi2196 & w5326;
assign w7736 = ~w7734 & ~w7735;
assign w7737 = pi1801 & ~w5100;
assign w7738 = pi2195 & w5100;
assign w7739 = ~w7737 & ~w7738;
assign w7740 = pi1802 & ~w6718;
assign w7741 = pi2172 & w6718;
assign w7742 = ~w7740 & ~w7741;
assign w7743 = pi1803 & ~w5100;
assign w7744 = pi2167 & w5100;
assign w7745 = ~w7743 & ~w7744;
assign w7746 = pi1804 & ~w5326;
assign w7747 = pi2191 & w5326;
assign w7748 = ~w7746 & ~w7747;
assign w7749 = pi1805 & ~w6567;
assign w7750 = pi2195 & w6567;
assign w7751 = ~w7749 & ~w7750;
assign w7752 = pi1806 & ~w5190;
assign w7753 = pi2171 & w5190;
assign w7754 = ~w7752 & ~w7753;
assign w7755 = pi1807 & ~w5315;
assign w7756 = pi2171 & w5315;
assign w7757 = ~w7755 & ~w7756;
assign w7758 = pi1808 & ~w5190;
assign w7759 = pi2193 & w5190;
assign w7760 = ~w7758 & ~w7759;
assign w7761 = pi1809 & ~w5100;
assign w7762 = pi2179 & w5100;
assign w7763 = ~w7761 & ~w7762;
assign w7764 = pi1810 & ~w5100;
assign w7765 = pi2170 & w5100;
assign w7766 = ~w7764 & ~w7765;
assign w7767 = pi1811 & ~w5100;
assign w7768 = pi2191 & w5100;
assign w7769 = ~w7767 & ~w7768;
assign w7770 = pi1812 & ~w5100;
assign w7771 = pi2176 & w5100;
assign w7772 = ~w7770 & ~w7771;
assign w7773 = pi1813 & ~w5100;
assign w7774 = pi2178 & w5100;
assign w7775 = ~w7773 & ~w7774;
assign w7776 = pi1814 & ~w5326;
assign w7777 = pi2181 & w5326;
assign w7778 = ~w7776 & ~w7777;
assign w7779 = pi1815 & ~w5190;
assign w7780 = pi2185 & w5190;
assign w7781 = ~w7779 & ~w7780;
assign w7782 = pi1816 & ~w5100;
assign w7783 = pi2172 & w5100;
assign w7784 = ~w7782 & ~w7783;
assign w7785 = pi1817 & ~w6567;
assign w7786 = pi2191 & w6567;
assign w7787 = ~w7785 & ~w7786;
assign w7788 = pi1818 & ~w5190;
assign w7789 = pi2168 & w5190;
assign w7790 = ~w7788 & ~w7789;
assign w7791 = pi1819 & ~w6567;
assign w7792 = pi2170 & w6567;
assign w7793 = ~w7791 & ~w7792;
assign w7794 = pi1820 & ~w5326;
assign w7795 = pi2176 & w5326;
assign w7796 = ~w7794 & ~w7795;
assign w7797 = pi1821 & ~w5406;
assign w7798 = pi2178 & w5406;
assign w7799 = ~w7797 & ~w7798;
assign w7800 = pi1822 & ~w5402;
assign w7801 = pi2191 & w5402;
assign w7802 = ~w7800 & ~w7801;
assign w7803 = pi1823 & ~w6567;
assign w7804 = pi2172 & w6567;
assign w7805 = ~w7803 & ~w7804;
assign w7806 = pi1824 & ~w5422;
assign w7807 = pi2170 & w5422;
assign w7808 = ~w7806 & ~w7807;
assign w7809 = pi1825 & ~w6567;
assign w7810 = pi2179 & w6567;
assign w7811 = ~w7809 & ~w7810;
assign w7812 = pi1826 & ~w6567;
assign w7813 = pi2176 & w6567;
assign w7814 = ~w7812 & ~w7813;
assign w7815 = pi1827 & ~w6567;
assign w7816 = pi2178 & w6567;
assign w7817 = ~w7815 & ~w7816;
assign w7818 = pi1828 & ~w5385;
assign w7819 = pi2194 & w5385;
assign w7820 = ~w7818 & ~w7819;
assign w7821 = pi1829 & ~w5402;
assign w7822 = pi2195 & w5402;
assign w7823 = ~w7821 & ~w7822;
assign w7824 = pi1830 & ~w5402;
assign w7825 = pi2167 & w5402;
assign w7826 = ~w7824 & ~w7825;
assign w7827 = pi1831 & ~w5326;
assign w7828 = pi2198 & w5326;
assign w7829 = ~w7827 & ~w7828;
assign w7830 = ~pi1989 & w4937;
assign w7831 = pi1832 & ~w7830;
assign w7832 = pi2172 & w7830;
assign w7833 = ~w7831 & ~w7832;
assign w7834 = pi1833 & ~w5315;
assign w7835 = pi2186 & w5315;
assign w7836 = ~w7834 & ~w7835;
assign w7837 = pi1159 & w4931;
assign w7838 = pi1975 & w4918;
assign w7839 = pi2082 & w4939;
assign w7840 = w4924 & w4925;
assign w7841 = pi2119 & w7840;
assign w7842 = pi1131 & w4935;
assign w7843 = pi1873 & w4937;
assign w7844 = pi1210 & w4915;
assign w7845 = pi2151 & w4933;
assign w7846 = pi2050 & w4921;
assign w7847 = ~w7837 & ~w7842;
assign w7848 = ~w7843 & ~w7844;
assign w7849 = ~w7845 & w7848;
assign w7850 = ~w7838 & w7847;
assign w7851 = ~w7839 & ~w7841;
assign w7852 = ~w7846 & w7851;
assign w7853 = w7849 & w7850;
assign w7854 = w7852 & w7853;
assign w7855 = pi1848 & w4937;
assign w7856 = pi1977 & w4918;
assign w7857 = pi2121 & w7840;
assign w7858 = pi2084 & w4939;
assign w7859 = pi1185 & w4935;
assign w7860 = pi1161 & w4931;
assign w7861 = pi2143 & w4933;
assign w7862 = pi1208 & w4915;
assign w7863 = pi2051 & w4921;
assign w7864 = ~w7855 & ~w7859;
assign w7865 = ~w7860 & ~w7861;
assign w7866 = ~w7862 & w7865;
assign w7867 = ~w7856 & w7864;
assign w7868 = ~w7857 & ~w7858;
assign w7869 = ~w7863 & w7868;
assign w7870 = w7866 & w7867;
assign w7871 = w7869 & w7870;
assign w7872 = pi1165 & w4935;
assign w7873 = pi1964 & w4918;
assign w7874 = pi2129 & w4939;
assign w7875 = pi2092 & w7840;
assign w7876 = pi1189 & w4915;
assign w7877 = pi2149 & w4933;
assign w7878 = pi1840 & w4937;
assign w7879 = pi1146 & w4931;
assign w7880 = pi2040 & w4921;
assign w7881 = ~w7872 & ~w7876;
assign w7882 = ~w7877 & ~w7878;
assign w7883 = ~w7879 & w7882;
assign w7884 = ~w7873 & w7881;
assign w7885 = ~w7874 & ~w7875;
assign w7886 = ~w7880 & w7885;
assign w7887 = w7883 & w7884;
assign w7888 = w7886 & w7887;
assign w7889 = pi1838 & ~w7830;
assign w7890 = pi2195 & w7830;
assign w7891 = ~w7889 & ~w7890;
assign w7892 = pi1839 & ~w7830;
assign w7893 = pi2186 & w7830;
assign w7894 = ~w7892 & ~w7893;
assign w7895 = pi1840 & ~w7830;
assign w7896 = pi2183 & w7830;
assign w7897 = ~w7895 & ~w7896;
assign w7898 = pi1841 & ~w7830;
assign w7899 = pi2168 & w7830;
assign w7900 = ~w7898 & ~w7899;
assign w7901 = pi1842 & ~w7830;
assign w7902 = pi2174 & w7830;
assign w7903 = ~w7901 & ~w7902;
assign w7904 = pi1843 & ~w7830;
assign w7905 = pi2197 & w7830;
assign w7906 = ~w7904 & ~w7905;
assign w7907 = pi1844 & ~w7830;
assign w7908 = pi2198 & w7830;
assign w7909 = ~w7907 & ~w7908;
assign w7910 = pi1845 & ~w7830;
assign w7911 = pi2191 & w7830;
assign w7912 = ~w7910 & ~w7911;
assign w7913 = pi1846 & ~w7830;
assign w7914 = pi2194 & w7830;
assign w7915 = ~w7913 & ~w7914;
assign w7916 = pi1847 & ~w7830;
assign w7917 = pi2188 & w7830;
assign w7918 = ~w7916 & ~w7917;
assign w7919 = pi1848 & ~w7830;
assign w7920 = pi2184 & w7830;
assign w7921 = ~w7919 & ~w7920;
assign w7922 = pi1849 & ~w7830;
assign w7923 = pi2166 & w7830;
assign w7924 = ~w7922 & ~w7923;
assign w7925 = pi1850 & pi2035;
assign w7926 = pi1928 & ~pi2035;
assign w7927 = ~w7925 & ~w7926;
assign w7928 = pi1851 & pi2056;
assign w7929 = pi1928 & ~pi2056;
assign w7930 = ~w7928 & ~w7929;
assign w7931 = pi1852 & pi2057;
assign w7932 = pi1928 & ~pi2057;
assign w7933 = ~w7931 & ~w7932;
assign w7934 = pi1853 & pi2059;
assign w7935 = pi1928 & ~pi2059;
assign w7936 = ~w7934 & ~w7935;
assign w7937 = pi1854 & ~w5315;
assign w7938 = pi2197 & w5315;
assign w7939 = ~w7937 & ~w7938;
assign w7940 = pi1855 & ~w5315;
assign w7941 = pi2166 & w5315;
assign w7942 = ~w7940 & ~w7941;
assign w7943 = pi1931 & pi2033;
assign w7944 = pi1856 & ~pi1931;
assign w7945 = ~w7943 & ~w7944;
assign w7946 = pi1857 & pi1943;
assign w7947 = ~pi1943 & pi2020;
assign w7948 = ~w7946 & ~w7947;
assign w7949 = pi1188 & w4915;
assign w7950 = pi1948 & w4918;
assign w7951 = pi2127 & w4939;
assign w7952 = pi2039 & w4921;
assign w7953 = pi2156 & w4933;
assign w7954 = pi1164 & w4935;
assign w7955 = pi1145 & w4931;
assign w7956 = pi1839 & w4937;
assign w7957 = pi2091 & w7840;
assign w7958 = ~w7949 & ~w7953;
assign w7959 = ~w7954 & ~w7955;
assign w7960 = ~w7956 & w7959;
assign w7961 = ~w7950 & w7958;
assign w7962 = ~w7951 & ~w7952;
assign w7963 = ~w7957 & w7962;
assign w7964 = w7960 & w7961;
assign w7965 = w7963 & w7964;
assign w7966 = pi2148 & w4933;
assign w7967 = pi0248 & w4918;
assign w7968 = pi2062 & w4939;
assign w7969 = pi2021 & w4921;
assign w7970 = pi1193 & w4915;
assign w7971 = pi1168 & w4935;
assign w7972 = pi1843 & w4937;
assign w7973 = pi1149 & w4931;
assign w7974 = pi2097 & w7840;
assign w7975 = ~w7966 & ~w7970;
assign w7976 = ~w7971 & ~w7972;
assign w7977 = ~w7973 & w7976;
assign w7978 = ~w7967 & w7975;
assign w7979 = ~w7968 & ~w7969;
assign w7980 = ~w7974 & w7979;
assign w7981 = w7977 & w7978;
assign w7982 = w7980 & w7981;
assign w7983 = pi2154 & w4933;
assign w7984 = pi1966 & w4918;
assign w7985 = pi2095 & w7840;
assign w7986 = pi2042 & w4921;
assign w7987 = pi1842 & w4937;
assign w7988 = pi1167 & w4935;
assign w7989 = pi1148 & w4931;
assign w7990 = pi1192 & w4915;
assign w7991 = pi2090 & w4939;
assign w7992 = ~w7983 & ~w7987;
assign w7993 = ~w7988 & ~w7989;
assign w7994 = ~w7990 & w7993;
assign w7995 = ~w7984 & w7992;
assign w7996 = ~w7985 & ~w7986;
assign w7997 = ~w7991 & w7996;
assign w7998 = w7994 & w7995;
assign w7999 = w7997 & w7998;
assign w8000 = pi1147 & w4931;
assign w8001 = pi1965 & w4918;
assign w8002 = pi2128 & w4939;
assign w8003 = pi2041 & w4921;
assign w8004 = pi1841 & w4937;
assign w8005 = pi1166 & w4935;
assign w8006 = pi2145 & w4933;
assign w8007 = pi1191 & w4915;
assign w8008 = pi2094 & w7840;
assign w8009 = ~w8000 & ~w8004;
assign w8010 = ~w8005 & ~w8006;
assign w8011 = ~w8007 & w8010;
assign w8012 = ~w8001 & w8009;
assign w8013 = ~w8002 & ~w8003;
assign w8014 = ~w8008 & w8013;
assign w8015 = w8011 & w8012;
assign w8016 = w8014 & w8015;
assign w8017 = pi1832 & w4937;
assign w8018 = pi0229 & w4918;
assign w8019 = pi2038 & w4921;
assign w8020 = pi2061 & w4939;
assign w8021 = pi2153 & w4933;
assign w8022 = pi1020 & w4935;
assign w8023 = pi1134 & w4931;
assign w8024 = pi1190 & w4915;
assign w8025 = pi2093 & w7840;
assign w8026 = ~w8017 & ~w8021;
assign w8027 = ~w8022 & ~w8023;
assign w8028 = ~w8024 & w8027;
assign w8029 = ~w8018 & w8026;
assign w8030 = ~w8019 & ~w8020;
assign w8031 = ~w8025 & w8030;
assign w8032 = w8028 & w8029;
assign w8033 = w8031 & w8032;
assign w8034 = pi2144 & w4933;
assign w8035 = pi1982 & w4918;
assign w8036 = pi2087 & w4939;
assign w8037 = pi2124 & w7840;
assign w8038 = pi1187 & w4935;
assign w8039 = pi1209 & w4915;
assign w8040 = pi1163 & w4931;
assign w8041 = pi1870 & w4937;
assign w8042 = pi2054 & w4921;
assign w8043 = ~w8034 & ~w8038;
assign w8044 = ~w8039 & ~w8040;
assign w8045 = ~w8041 & w8044;
assign w8046 = ~w8035 & w8043;
assign w8047 = ~w8036 & ~w8037;
assign w8048 = ~w8042 & w8047;
assign w8049 = w8045 & w8046;
assign w8050 = w8048 & w8049;
assign w8051 = pi1186 & w4935;
assign w8052 = pi1976 & w4918;
assign w8053 = pi2122 & w7840;
assign w8054 = pi2085 & w4939;
assign w8055 = pi2147 & w4933;
assign w8056 = pi1132 & w4915;
assign w8057 = pi1849 & w4937;
assign w8058 = pi1162 & w4931;
assign w8059 = pi2052 & w4921;
assign w8060 = ~w8051 & ~w8055;
assign w8061 = ~w8056 & ~w8057;
assign w8062 = ~w8058 & w8061;
assign w8063 = ~w8052 & w8060;
assign w8064 = ~w8053 & ~w8054;
assign w8065 = ~w8059 & w8064;
assign w8066 = w8062 & w8063;
assign w8067 = w8065 & w8066;
assign w8068 = pi1137 & w4931;
assign w8069 = pi1950 & w4918;
assign w8070 = pi2098 & w7840;
assign w8071 = pi2125 & w4939;
assign w8072 = pi1211 & w4915;
assign w8073 = pi1821 & w4935;
assign w8074 = pi2150 & w4933;
assign w8075 = pi1871 & w4937;
assign w8076 = pi2022 & w4921;
assign w8077 = ~w8068 & ~w8072;
assign w8078 = ~w8073 & ~w8074;
assign w8079 = ~w8075 & w8078;
assign w8080 = ~w8069 & w8077;
assign w8081 = ~w8070 & ~w8071;
assign w8082 = ~w8076 & w8081;
assign w8083 = w8079 & w8080;
assign w8084 = w8082 & w8083;
assign w8085 = pi1160 & w4931;
assign w8086 = pi0230 & w4918;
assign w8087 = pi2120 & w7840;
assign w8088 = pi2083 & w4939;
assign w8089 = pi1184 & w4935;
assign w8090 = pi1207 & w4915;
assign w8091 = pi1847 & w4937;
assign w8092 = pi2157 & w4933;
assign w8093 = pi2103 & w4921;
assign w8094 = ~w8085 & ~w8089;
assign w8095 = ~w8090 & ~w8091;
assign w8096 = ~w8092 & w8095;
assign w8097 = ~w8086 & w8094;
assign w8098 = ~w8087 & ~w8088;
assign w8099 = ~w8093 & w8098;
assign w8100 = w8096 & w8097;
assign w8101 = w8099 & w8100;
assign w8102 = pi1779 & w4915;
assign w8103 = pi1974 & w4918;
assign w8104 = pi2049 & w4921;
assign w8105 = pi2118 & w7840;
assign w8106 = pi1183 & w4935;
assign w8107 = pi1846 & w4937;
assign w8108 = pi1158 & w4931;
assign w8109 = pi2160 & w4933;
assign w8110 = pi2080 & w4939;
assign w8111 = ~w8102 & ~w8106;
assign w8112 = ~w8107 & ~w8108;
assign w8113 = ~w8109 & w8112;
assign w8114 = ~w8103 & w8111;
assign w8115 = ~w8104 & ~w8105;
assign w8116 = ~w8110 & w8115;
assign w8117 = w8113 & w8114;
assign w8118 = w8116 & w8117;
assign w8119 = pi1036 & w4931;
assign w8120 = pi0251 & w4918;
assign w8121 = pi2123 & w7840;
assign w8122 = pi2086 & w4939;
assign w8123 = pi1838 & w4937;
assign w8124 = pi1690 & w4915;
assign w8125 = pi1035 & w4935;
assign w8126 = pi2152 & w4933;
assign w8127 = pi2053 & w4921;
assign w8128 = ~w8119 & ~w8123;
assign w8129 = ~w8124 & ~w8125;
assign w8130 = ~w8126 & w8129;
assign w8131 = ~w8120 & w8128;
assign w8132 = ~w8121 & ~w8122;
assign w8133 = ~w8127 & w8132;
assign w8134 = w8130 & w8131;
assign w8135 = w8133 & w8134;
assign w8136 = pi1206 & w4915;
assign w8137 = pi0250 & w4918;
assign w8138 = pi2115 & w7840;
assign w8139 = pi2047 & w4921;
assign w8140 = pi2155 & w4933;
assign w8141 = pi1157 & w4931;
assign w8142 = pi1845 & w4937;
assign w8143 = pi1130 & w4935;
assign w8144 = pi2077 & w4939;
assign w8145 = ~w8136 & ~w8140;
assign w8146 = ~w8141 & ~w8142;
assign w8147 = ~w8143 & w8146;
assign w8148 = ~w8137 & w8145;
assign w8149 = ~w8138 & ~w8139;
assign w8150 = ~w8144 & w8149;
assign w8151 = w8147 & w8148;
assign w8152 = w8150 & w8151;
assign w8153 = pi1870 & ~w7830;
assign w8154 = pi2192 & w7830;
assign w8155 = ~w8153 & ~w8154;
assign w8156 = pi1871 & ~w7830;
assign w8157 = pi2178 & w7830;
assign w8158 = ~w8156 & ~w8157;
assign w8159 = pi1872 & ~w5315;
assign w8160 = pi2173 & w5315;
assign w8161 = ~w8159 & ~w8160;
assign w8162 = pi1873 & ~w7830;
assign w8163 = pi2167 & w7830;
assign w8164 = ~w8162 & ~w8163;
assign w8165 = pi1929 & pi2032;
assign w8166 = ~pi0259 & ~pi2032;
assign w8167 = ~w8165 & ~w8166;
assign w8168 = pi1875 & pi2058;
assign w8169 = pi1928 & ~pi2058;
assign w8170 = ~w8168 & ~w8169;
assign w8171 = pi1877 & pi1952;
assign w8172 = ~pi1952 & pi2055;
assign w8173 = ~w8171 & ~w8172;
assign w8174 = ~pi1989 & w4924;
assign w8175 = pi2186 & w8174;
assign w8176 = pi2198 & w8174;
assign w8177 = pi1144 & w4933;
assign w8178 = pi1182 & w4935;
assign w8179 = pi2117 & w7840;
assign w8180 = pi2096 & w4921;
assign w8181 = pi2079 & w4939;
assign w8182 = ~w8177 & ~w8178;
assign w8183 = ~w8179 & w8182;
assign w8184 = ~w8180 & ~w8181;
assign w8185 = w8183 & w8184;
assign w8186 = pi1883 & pi2059;
assign w8187 = pi1942 & ~pi2059;
assign w8188 = ~w8186 & ~w8187;
assign w8189 = pi1884 & pi2035;
assign w8190 = pi1942 & ~pi2035;
assign w8191 = ~w8189 & ~w8190;
assign w8192 = pi1885 & pi2056;
assign w8193 = pi1942 & ~pi2056;
assign w8194 = ~w8192 & ~w8193;
assign w8195 = pi1886 & pi2057;
assign w8196 = pi1942 & ~pi2057;
assign w8197 = ~w8195 & ~w8196;
assign w8198 = pi1201 & w4915;
assign w8199 = pi1156 & w4931;
assign w8200 = pi1175 & w4935;
assign w8201 = pi2030 & w4921;
assign w8202 = pi0841 & w4918;
assign w8203 = pi2068 & w4939;
assign w8204 = pi2108 & w7840;
assign w8205 = ~w8198 & ~w8199;
assign w8206 = ~w8200 & w8205;
assign w8207 = ~w8201 & ~w8202;
assign w8208 = ~w8203 & ~w8204;
assign w8209 = w8207 & w8208;
assign w8210 = w8206 & w8209;
assign w8211 = pi1970 & w4918;
assign w8212 = pi1133 & w4915;
assign w8213 = pi1012 & w4933;
assign w8214 = pi1762 & w4935;
assign w8215 = pi1128 & w4931;
assign w8216 = pi2029 & w4921;
assign w8217 = pi2067 & w4939;
assign w8218 = pi2107 & w7840;
assign w8219 = ~w8212 & ~w8213;
assign w8220 = ~w8214 & ~w8215;
assign w8221 = w8219 & w8220;
assign w8222 = ~w8211 & ~w8216;
assign w8223 = ~w8217 & ~w8218;
assign w8224 = w8222 & w8223;
assign w8225 = w8221 & w8224;
assign w8226 = pi1946 & w4918;
assign w8227 = pi1174 & w4935;
assign w8228 = pi1155 & w4931;
assign w8229 = pi1200 & w4915;
assign w8230 = pi1143 & w4933;
assign w8231 = pi2028 & w4921;
assign w8232 = pi2106 & w7840;
assign w8233 = pi2066 & w4939;
assign w8234 = ~w8227 & ~w8228;
assign w8235 = ~w8229 & ~w8230;
assign w8236 = w8234 & w8235;
assign w8237 = ~w8226 & ~w8231;
assign w8238 = ~w8232 & ~w8233;
assign w8239 = w8237 & w8238;
assign w8240 = w8236 & w8239;
assign w8241 = pi1967 & w4918;
assign w8242 = pi1194 & w4915;
assign w8243 = pi1139 & w4933;
assign w8244 = pi1169 & w4935;
assign w8245 = pi1150 & w4931;
assign w8246 = pi2099 & w7840;
assign w8247 = pi2072 & w4921;
assign w8248 = pi2071 & w4939;
assign w8249 = ~w8242 & ~w8243;
assign w8250 = ~w8244 & ~w8245;
assign w8251 = w8249 & w8250;
assign w8252 = ~w8241 & ~w8246;
assign w8253 = ~w8247 & ~w8248;
assign w8254 = w8252 & w8253;
assign w8255 = w8251 & w8254;
assign w8256 = pi0842 & w4918;
assign w8257 = pi1173 & w4935;
assign w8258 = pi1142 & w4933;
assign w8259 = pi1154 & w4931;
assign w8260 = pi1199 & w4915;
assign w8261 = pi2027 & w4921;
assign w8262 = pi2105 & w7840;
assign w8263 = pi2065 & w4939;
assign w8264 = ~w8257 & ~w8258;
assign w8265 = ~w8259 & ~w8260;
assign w8266 = w8264 & w8265;
assign w8267 = ~w8256 & ~w8261;
assign w8268 = ~w8262 & ~w8263;
assign w8269 = w8267 & w8268;
assign w8270 = w8266 & w8269;
assign w8271 = pi1969 & w4918;
assign w8272 = pi1138 & w4931;
assign w8273 = pi1141 & w4933;
assign w8274 = pi1197 & w4915;
assign w8275 = pi1789 & w4935;
assign w8276 = pi2064 & w4939;
assign w8277 = pi2025 & w4921;
assign w8278 = pi2102 & w7840;
assign w8279 = ~w8272 & ~w8273;
assign w8280 = ~w8274 & ~w8275;
assign w8281 = w8279 & w8280;
assign w8282 = ~w8271 & ~w8276;
assign w8283 = ~w8277 & ~w8278;
assign w8284 = w8282 & w8283;
assign w8285 = w8281 & w8284;
assign w8286 = pi0249 & w4918;
assign w8287 = pi1151 & w4931;
assign w8288 = pi1170 & w4935;
assign w8289 = pi1140 & w4933;
assign w8290 = pi1195 & w4915;
assign w8291 = pi2023 & w4921;
assign w8292 = pi2126 & w4939;
assign w8293 = pi2100 & w7840;
assign w8294 = ~w8287 & ~w8288;
assign w8295 = ~w8289 & ~w8290;
assign w8296 = w8294 & w8295;
assign w8297 = ~w8286 & ~w8291;
assign w8298 = ~w8292 & ~w8293;
assign w8299 = w8297 & w8298;
assign w8300 = w8296 & w8299;
assign w8301 = pi1971 & w4918;
assign w8302 = pi1176 & w4935;
assign w8303 = pi1202 & w4915;
assign w8304 = pi2109 & w7840;
assign w8305 = pi2069 & w4939;
assign w8306 = pi2088 & w4921;
assign w8307 = ~w8302 & ~w8303;
assign w8308 = ~w8301 & w8307;
assign w8309 = ~w8304 & ~w8305;
assign w8310 = ~w8306 & w8309;
assign w8311 = w8308 & w8310;
assign w8312 = pi1181 & w4935;
assign w8313 = pi2078 & w4939;
assign w8314 = pi2048 & w4921;
assign w8315 = pi2116 & w7840;
assign w8316 = ~w8312 & ~w8313;
assign w8317 = ~w8314 & ~w8315;
assign w8318 = w8316 & w8317;
assign w8319 = pi1973 & w4918;
assign w8320 = pi1205 & w4915;
assign w8321 = pi1179 & w4935;
assign w8322 = pi2075 & w4939;
assign w8323 = pi2045 & w4921;
assign w8324 = pi2113 & w7840;
assign w8325 = ~w8320 & ~w8321;
assign w8326 = ~w8319 & w8325;
assign w8327 = ~w8322 & ~w8323;
assign w8328 = ~w8324 & w8327;
assign w8329 = w8326 & w8328;
assign w8330 = pi1949 & w4918;
assign w8331 = pi1204 & w4915;
assign w8332 = pi1178 & w4935;
assign w8333 = pi2044 & w4921;
assign w8334 = pi2112 & w7840;
assign w8335 = pi2074 & w4939;
assign w8336 = ~w8331 & ~w8332;
assign w8337 = ~w8330 & w8336;
assign w8338 = ~w8333 & ~w8334;
assign w8339 = ~w8335 & w8338;
assign w8340 = w8337 & w8339;
assign w8341 = pi0815 & w4918;
assign w8342 = pi1760 & w4915;
assign w8343 = pi1777 & w4935;
assign w8344 = pi2073 & w4939;
assign w8345 = pi2111 & w7840;
assign w8346 = pi2089 & w4921;
assign w8347 = ~w8342 & ~w8343;
assign w8348 = ~w8341 & w8347;
assign w8349 = ~w8344 & ~w8345;
assign w8350 = ~w8346 & w8349;
assign w8351 = w8348 & w8350;
assign w8352 = pi1180 & w4935;
assign w8353 = pi2076 & w4939;
assign w8354 = pi2114 & w7840;
assign w8355 = pi2046 & w4921;
assign w8356 = ~w8352 & ~w8353;
assign w8357 = ~w8354 & ~w8355;
assign w8358 = w8356 & w8357;
assign w8359 = pi1972 & w4918;
assign w8360 = pi1177 & w4935;
assign w8361 = pi1203 & w4915;
assign w8362 = pi2070 & w4939;
assign w8363 = pi2043 & w4921;
assign w8364 = pi2110 & w7840;
assign w8365 = ~w8360 & ~w8361;
assign w8366 = ~w8359 & w8365;
assign w8367 = ~w8362 & ~w8363;
assign w8368 = ~w8364 & w8367;
assign w8369 = w8366 & w8368;
assign w8370 = pi1901 & pi2058;
assign w8371 = pi1942 & ~pi2058;
assign w8372 = ~w8370 & ~w8371;
assign w8373 = pi1968 & w4918;
assign w8374 = pi1171 & w4935;
assign w8375 = pi1771 & w4933;
assign w8376 = pi1196 & w4915;
assign w8377 = pi1152 & w4931;
assign w8378 = pi2024 & w4921;
assign w8379 = pi2063 & w4939;
assign w8380 = pi2101 & w7840;
assign w8381 = ~w8374 & ~w8375;
assign w8382 = ~w8376 & ~w8377;
assign w8383 = w8381 & w8382;
assign w8384 = ~w8373 & ~w8378;
assign w8385 = ~w8379 & ~w8380;
assign w8386 = w8384 & w8385;
assign w8387 = w8383 & w8386;
assign w8388 = ~w4961 & w4966;
assign w8389 = pi0353 & w8388;
assign w8390 = ~w4962 & ~w4966;
assign w8391 = pi0353 & ~w604;
assign w8392 = ~w4963 & ~w8391;
assign w8393 = pi0353 & w2282;
assign w8394 = w4969 & ~w8393;
assign w8395 = ~w4969 & w8393;
assign w8396 = ~w8394 & ~w8395;
assign w8397 = ~w8390 & ~w8392;
assign w8398 = ~w8389 & w8397;
assign w8399 = ~w8396 & w8398;
assign w8400 = ~w4988 & ~w4992;
assign w8401 = w725 & w4995;
assign w8402 = ~w4987 & w4992;
assign w8403 = ~w639 & ~w8401;
assign w8404 = ~w8402 & w8403;
assign w8405 = pi0262 & ~w8404;
assign w8406 = w4989 & w4995;
assign w8407 = ~pi0262 & ~w8406;
assign w8408 = ~w725 & ~w4995;
assign w8409 = ~w8400 & ~w8408;
assign w8410 = ~w8407 & w8409;
assign w8411 = ~w8405 & w8410;
assign w8412 = ~w4951 & ~w4955;
assign w8413 = w813 & w4950;
assign w8414 = ~w631 & ~w4956;
assign w8415 = ~w8413 & w8414;
assign w8416 = pi0261 & ~w8415;
assign w8417 = ~w4951 & ~w4952;
assign w8418 = w4950 & w8417;
assign w8419 = ~pi0261 & ~w8418;
assign w8420 = ~w813 & ~w4950;
assign w8421 = ~w8412 & ~w8420;
assign w8422 = ~w8419 & w8421;
assign w8423 = ~w8416 & w8422;
assign w8424 = ~w5018 & ~w5022;
assign w8425 = w714 & w5017;
assign w8426 = ~w611 & ~w5023;
assign w8427 = ~w8425 & w8426;
assign w8428 = pi0354 & ~w8427;
assign w8429 = ~pi0354 & ~w5024;
assign w8430 = pi0354 & w714;
assign w8431 = ~w5017 & ~w8430;
assign w8432 = ~w8424 & ~w8431;
assign w8433 = ~w8429 & w8432;
assign w8434 = ~w8428 & w8433;
assign w8435 = ~w4975 & ~w4979;
assign w8436 = w773 & w4982;
assign w8437 = ~w4974 & w4979;
assign w8438 = ~w647 & ~w8436;
assign w8439 = ~w8437 & w8438;
assign w8440 = pi0263 & ~w8439;
assign w8441 = w4976 & w4982;
assign w8442 = ~pi0263 & ~w8441;
assign w8443 = ~w773 & ~w4982;
assign w8444 = ~w8435 & ~w8443;
assign w8445 = ~w8442 & w8444;
assign w8446 = ~w8440 & w8445;
assign w8447 = ~w5007 & ~w5008;
assign w8448 = w5004 & w5011;
assign w8449 = ~pi0260 & ~w8448;
assign w8450 = ~w863 & ~w5004;
assign w8451 = w5007 & ~w5009;
assign w8452 = w863 & w5004;
assign w8453 = ~w623 & ~w8451;
assign w8454 = ~w8452 & w8453;
assign w8455 = pi0260 & ~w8454;
assign w8456 = ~w8447 & ~w8450;
assign w8457 = ~w8449 & w8456;
assign w8458 = ~w8455 & w8457;
assign w8459 = pi1917 & pi1921;
assign w8460 = ~pi2031 & w8459;
assign w8461 = ~pi1911 & ~w8460;
assign w8462 = pi1911 & w8460;
assign w8463 = pi1036 & ~w8461;
assign w8464 = ~w8462 & w8463;
assign w8465 = pi1915 & pi1918;
assign w8466 = ~pi2034 & w8465;
assign w8467 = ~pi1912 & ~w8466;
assign w8468 = pi1912 & w8466;
assign w8469 = pi1150 & ~w8467;
assign w8470 = ~w8468 & w8469;
assign w8471 = ~pi2010 & ~pi2036;
assign w8472 = ~pi1913 & ~w8471;
assign w8473 = ~pi2009 & ~pi2031;
assign w8474 = ~pi1914 & ~w8473;
assign w8475 = pi1918 & ~pi2034;
assign w8476 = ~pi1915 & ~w8475;
assign w8477 = pi1150 & ~w8466;
assign w8478 = ~w8476 & w8477;
assign w8479 = pi1916 & pi1919;
assign w8480 = ~pi2036 & w8479;
assign w8481 = pi1919 & ~pi2036;
assign w8482 = ~pi1916 & ~w8481;
assign w8483 = pi1145 & ~w8480;
assign w8484 = ~w8482 & w8483;
assign w8485 = pi1921 & ~pi2031;
assign w8486 = ~pi1917 & ~w8485;
assign w8487 = pi1036 & ~w8460;
assign w8488 = ~w8486 & w8487;
assign w8489 = ~pi1918 & pi2034;
assign w8490 = pi1150 & ~w8475;
assign w8491 = ~w8489 & w8490;
assign w8492 = ~pi1919 & pi2036;
assign w8493 = pi1145 & ~w8481;
assign w8494 = ~w8492 & w8493;
assign w8495 = ~pi1920 & ~w8480;
assign w8496 = pi1920 & w8480;
assign w8497 = pi1145 & ~w8495;
assign w8498 = ~w8496 & w8497;
assign w8499 = ~pi1921 & pi2031;
assign w8500 = pi1036 & ~w8485;
assign w8501 = ~w8499 & w8500;
assign w8502 = pi1922 & pi2035;
assign w8503 = pi1992 & ~pi2035;
assign w8504 = ~w8502 & ~w8503;
assign w8505 = pi1923 & pi2056;
assign w8506 = pi1992 & ~pi2056;
assign w8507 = ~w8505 & ~w8506;
assign w8508 = pi1924 & pi2057;
assign w8509 = pi1992 & ~pi2057;
assign w8510 = ~w8508 & ~w8509;
assign w8511 = pi1925 & pi2059;
assign w8512 = pi1992 & ~pi2059;
assign w8513 = ~w8511 & ~w8512;
assign w8514 = pi1926 & pi2058;
assign w8515 = pi1992 & ~pi2058;
assign w8516 = ~w8514 & ~w8515;
assign w8517 = ~pi2018 & ~pi2034;
assign w8518 = ~pi1927 & ~w8517;
assign w8519 = ~pi0257 & ~pi2032;
assign w8520 = pi1932 & pi2056;
assign w8521 = pi2014 & ~pi2056;
assign w8522 = ~w8520 & ~w8521;
assign w8523 = pi1933 & pi2059;
assign w8524 = pi2014 & ~pi2059;
assign w8525 = ~w8523 & ~w8524;
assign w8526 = pi1934 & pi2057;
assign w8527 = pi2014 & ~pi2057;
assign w8528 = ~w8526 & ~w8527;
assign w8529 = pi1935 & pi2058;
assign w8530 = pi2014 & ~pi2058;
assign w8531 = ~w8529 & ~w8530;
assign w8532 = pi2201 & w681;
assign w8533 = pi2013 & w8532;
assign w8534 = pi2162 & w8533;
assign w8535 = w4917 & w8534;
assign w8536 = w4931 & w8535;
assign w8537 = w4924 & w8535;
assign w8538 = w4935 & w8535;
assign w8539 = w4937 & w8535;
assign w8540 = w4933 & w8535;
assign w8541 = w4915 & w8535;
assign w8542 = pi1995 & pi1996;
assign w8543 = pi1986 & w8542;
assign w8544 = pi1955 & w8543;
assign w8545 = pi1957 & w8544;
assign w8546 = ~pi1944 & ~w8545;
assign w8547 = pi1944 & w8545;
assign w8548 = ~pi2133 & ~w8546;
assign w8549 = ~w8547 & w8548;
assign w8550 = pi0229 & pi1190;
assign w8551 = pi1192 & pi1966;
assign w8552 = pi1191 & pi1965;
assign w8553 = pi0842 & pi1199;
assign w8554 = pi0230 & pi1207;
assign w8555 = pi0251 & pi1690;
assign w8556 = pi1204 & pi1949;
assign w8557 = pi1202 & pi1971;
assign w8558 = pi1208 & pi1977;
assign w8559 = pi1210 & pi1975;
assign w8560 = pi1209 & pi1982;
assign w8561 = pi1133 & pi1970;
assign w8562 = pi1194 & pi1967;
assign w8563 = pi0248 & pi1193;
assign w8564 = pi1196 & pi1968;
assign w8565 = pi1189 & pi1964;
assign w8566 = pi1197 & pi1969;
assign w8567 = pi1779 & pi1974;
assign w8568 = pi1188 & pi1948;
assign w8569 = pi1200 & pi1946;
assign w8570 = pi1205 & pi1973;
assign w8571 = pi1132 & pi1976;
assign w8572 = pi0815 & pi1760;
assign w8573 = pi0841 & pi1201;
assign w8574 = pi1203 & pi1972;
assign w8575 = pi0810 & pi1198;
assign w8576 = pi0250 & pi1206;
assign w8577 = pi0249 & pi1195;
assign w8578 = pi1211 & pi1950;
assign w8579 = ~w8550 & ~w8551;
assign w8580 = ~w8552 & ~w8553;
assign w8581 = ~w8554 & ~w8555;
assign w8582 = ~w8556 & ~w8557;
assign w8583 = ~w8558 & ~w8559;
assign w8584 = ~w8560 & ~w8561;
assign w8585 = ~w8562 & ~w8563;
assign w8586 = ~w8564 & ~w8565;
assign w8587 = ~w8566 & ~w8567;
assign w8588 = ~w8568 & ~w8569;
assign w8589 = ~w8570 & ~w8571;
assign w8590 = ~w8572 & ~w8573;
assign w8591 = ~w8574 & ~w8575;
assign w8592 = ~w8576 & ~w8577;
assign w8593 = ~w8578 & w8592;
assign w8594 = w8590 & w8591;
assign w8595 = w8588 & w8589;
assign w8596 = w8586 & w8587;
assign w8597 = w8584 & w8585;
assign w8598 = w8582 & w8583;
assign w8599 = w8580 & w8581;
assign w8600 = w8579 & w8599;
assign w8601 = w8597 & w8598;
assign w8602 = w8595 & w8596;
assign w8603 = w8593 & w8594;
assign w8604 = w8602 & w8603;
assign w8605 = w8600 & w8601;
assign w8606 = w8604 & w8605;
assign w8607 = ~pi1913 & ~pi1946;
assign w8608 = ~w686 & ~w8607;
assign w8609 = pi1947 & pi2059;
assign w8610 = ~pi2059 & pi2164;
assign w8611 = ~w8609 & ~w8610;
assign w8612 = ~pi0873 & ~pi1948;
assign w8613 = ~w686 & ~w8612;
assign w8614 = ~pi1927 & ~pi1949;
assign w8615 = ~w686 & ~w8614;
assign w8616 = pi0452 & ~pi1950;
assign w8617 = ~w686 & ~w8616;
assign w8618 = pi1985 & pi1994;
assign w8619 = pi2000 & w8618;
assign w8620 = w8618 & w10744;
assign w8621 = pi1993 & w8620;
assign w8622 = pi1997 & w8621;
assign w8623 = ~pi1951 & pi1998;
assign w8624 = w8622 & w8623;
assign w8625 = pi1998 & w8622;
assign w8626 = pi1951 & ~w8625;
assign w8627 = ~pi2134 & ~w8624;
assign w8628 = ~w8626 & w8627;
assign w8629 = ~pi1955 & ~w8543;
assign w8630 = pi1995 & ~pi1996;
assign w8631 = pi1944 & ~pi1955;
assign w8632 = ~pi1957 & ~pi1986;
assign w8633 = w8631 & w8632;
assign w8634 = w8630 & w8633;
assign w8635 = ~pi2133 & ~w8634;
assign w8636 = ~w8544 & ~w8629;
assign w8637 = w8635 & w8636;
assign w8638 = w4890 & w10741;
assign w8639 = pi2003 & w8638;
assign w8640 = w8638 & w10742;
assign w8641 = ~pi1956 & ~w8640;
assign w8642 = pi1956 & w8640;
assign w8643 = pi0880 & ~w8641;
assign w8644 = ~w8642 & w8643;
assign w8645 = ~pi1957 & ~w8544;
assign w8646 = ~w8545 & w8635;
assign w8647 = ~w8645 & w8646;
assign w8648 = pi1958 & pi2059;
assign w8649 = ~pi2059 & pi2142;
assign w8650 = ~w8648 & ~w8649;
assign w8651 = pi1959 & pi2059;
assign w8652 = ~pi2059 & pi2161;
assign w8653 = ~w8651 & ~w8652;
assign w8654 = pi1960 & pi2057;
assign w8655 = ~pi2057 & pi2161;
assign w8656 = ~w8654 & ~w8655;
assign w8657 = pi1961 & pi2058;
assign w8658 = ~pi2058 & pi2161;
assign w8659 = ~w8657 & ~w8658;
assign w8660 = pi1962 & pi2058;
assign w8661 = ~pi2058 & pi2142;
assign w8662 = ~w8660 & ~w8661;
assign w8663 = ~w684 & ~w8534;
assign w8664 = ~pi1963 & ~w8663;
assign w8665 = pi0905 & ~pi1964;
assign w8666 = ~w686 & ~w8665;
assign w8667 = pi0451 & ~pi1965;
assign w8668 = ~w686 & ~w8667;
assign w8669 = pi0902 & ~pi1966;
assign w8670 = ~w686 & ~w8669;
assign w8671 = pi0901 & ~pi1967;
assign w8672 = ~w686 & ~w8671;
assign w8673 = pi0453 & ~pi1968;
assign w8674 = ~w686 & ~w8673;
assign w8675 = pi0904 & ~pi1969;
assign w8676 = ~w686 & ~w8675;
assign w8677 = pi0872 & ~pi1970;
assign w8678 = ~w686 & ~w8677;
assign w8679 = ~pi1914 & ~pi1971;
assign w8680 = ~w686 & ~w8679;
assign w8681 = pi0808 & ~pi1972;
assign w8682 = ~w686 & ~w8681;
assign w8683 = pi0636 & ~pi1973;
assign w8684 = ~w686 & ~w8683;
assign w8685 = pi0450 & ~pi1974;
assign w8686 = ~w686 & ~w8685;
assign w8687 = pi0899 & ~pi1975;
assign w8688 = ~w686 & ~w8687;
assign w8689 = pi0900 & ~pi1976;
assign w8690 = ~w686 & ~w8689;
assign w8691 = pi0806 & ~pi1977;
assign w8692 = ~w686 & ~w8691;
assign w8693 = pi1978 & pi2058;
assign w8694 = ~pi2058 & pi2081;
assign w8695 = ~w8693 & ~w8694;
assign w8696 = pi1979 & pi2058;
assign w8697 = ~pi2058 & pi2164;
assign w8698 = ~w8696 & ~w8697;
assign w8699 = pi1980 & pi2057;
assign w8700 = ~pi2057 & pi2081;
assign w8701 = ~w8699 & ~w8700;
assign w8702 = pi1981 & pi2059;
assign w8703 = ~pi2059 & pi2081;
assign w8704 = ~w8702 & ~w8703;
assign w8705 = pi0807 & ~pi1982;
assign w8706 = ~w686 & ~w8705;
assign w8707 = pi1983 & pi2057;
assign w8708 = ~pi2057 & pi2142;
assign w8709 = ~w8707 & ~w8708;
assign w8710 = pi1984 & pi2057;
assign w8711 = ~pi2057 & pi2164;
assign w8712 = ~w8710 & ~w8711;
assign w8713 = pi1985 & pi1999;
assign w8714 = ~pi1985 & ~pi1999;
assign w8715 = ~w8713 & ~w8714;
assign w8716 = ~pi2134 & ~w8715;
assign w8717 = ~pi1986 & ~w8542;
assign w8718 = ~w8543 & ~w8717;
assign w8719 = w8635 & w8718;
assign w8720 = w4961 & ~w4966;
assign w8721 = ~w8388 & ~w8720;
assign w8722 = w5019 & ~w5022;
assign w8723 = ~w5023 & ~w8722;
assign w8724 = w680 & w8534;
assign w8725 = ~pi1990 & ~w4891;
assign w8726 = pi0880 & ~w8638;
assign w8727 = ~w8725 & w8726;
assign w8728 = ~pi1993 & ~w8620;
assign w8729 = ~w8621 & ~w8728;
assign w8730 = ~pi2134 & ~w8729;
assign w8731 = pi2000 & w8713;
assign w8732 = ~pi1994 & ~w8731;
assign w8733 = ~w8620 & ~w8732;
assign w8734 = ~pi2134 & ~w8733;
assign w8735 = pi1995 & ~w8634;
assign w8736 = ~pi2133 & ~w8735;
assign w8737 = ~pi1995 & pi1996;
assign w8738 = ~w8630 & ~w8737;
assign w8739 = w8635 & ~w8738;
assign w8740 = ~pi1997 & ~w8621;
assign w8741 = ~w8622 & ~w8740;
assign w8742 = ~pi2134 & ~w8741;
assign w8743 = (~pi1998 & ~w8621) | (~pi1998 & w10743) | (~w8621 & w10743);
assign w8744 = ~w8625 & ~w8743;
assign w8745 = ~pi2134 & ~w8744;
assign w8746 = pi1999 & ~pi2134;
assign w8747 = ~pi2000 & ~w8713;
assign w8748 = ~w8731 & ~w8747;
assign w8749 = ~pi2134 & ~w8748;
assign w8750 = ~pi2001 & ~w8639;
assign w8751 = pi0880 & ~w8640;
assign w8752 = ~w8750 & w8751;
assign w8753 = ~pi1951 & ~pi1998;
assign w8754 = pi1994 & pi1997;
assign w8755 = ~pi1985 & ~pi2000;
assign w8756 = pi1993 & w8754;
assign w8757 = ~w8755 & w8756;
assign w8758 = w8753 & ~w8757;
assign w8759 = ~pi2003 & ~w8638;
assign w8760 = pi0880 & ~w8639;
assign w8761 = ~w8759 & w8760;
assign w8762 = w4952 & ~w4955;
assign w8763 = ~w4956 & ~w8762;
assign w8764 = w4987 & ~w4992;
assign w8765 = ~w8402 & ~w8764;
assign w8766 = w4974 & ~w4979;
assign w8767 = ~w8437 & ~w8766;
assign w8768 = ~w5007 & w5009;
assign w8769 = ~w8451 & ~w8768;
assign w8770 = ~pi0411 & pi1918;
assign w8771 = pi0412 & ~pi1915;
assign w8772 = ~pi0412 & pi1915;
assign w8773 = ~w8771 & ~w8772;
assign w8774 = w8770 & w8773;
assign w8775 = ~w8770 & ~w8773;
assign w8776 = ~w8774 & ~w8775;
assign w8777 = pi0463 & ~pi1911;
assign w8778 = ~pi0463 & pi1911;
assign w8779 = ~w8777 & ~w8778;
assign w8780 = pi0601 & ~pi1921;
assign w8781 = ~pi0601 & pi1921;
assign w8782 = ~w8780 & ~w8781;
assign w8783 = pi0602 & ~pi1917;
assign w8784 = ~pi0602 & pi1917;
assign w8785 = ~w8783 & ~w8784;
assign w8786 = w8782 & w8785;
assign w8787 = w3364 & w8779;
assign w8788 = w8786 & w8787;
assign w8789 = pi0643 & ~pi1920;
assign w8790 = ~pi0643 & pi1920;
assign w8791 = ~w8789 & ~w8790;
assign w8792 = pi0843 & ~pi1919;
assign w8793 = ~pi0843 & pi1919;
assign w8794 = ~w8792 & ~w8793;
assign w8795 = pi0746 & ~pi1916;
assign w8796 = ~pi0746 & pi1916;
assign w8797 = ~w8795 & ~w8796;
assign w8798 = w8794 & w8797;
assign w8799 = w3384 & w8791;
assign w8800 = w8798 & w8799;
assign w8801 = ~pi1993 & ~pi1997;
assign w8802 = ~pi1951 & w8801;
assign w8803 = ~w8619 & w8802;
assign w8804 = ~w8753 & ~w8803;
assign w8805 = ~pi2243 & ~pi2244;
assign w8806 = ~pi2245 & w8805;
assign w8807 = w8532 & w8806;
assign w8808 = ~w8534 & w8807;
assign w8809 = pi1994 & ~w8755;
assign w8810 = ~pi1998 & w8801;
assign w8811 = ~w8809 & w8810;
assign w8812 = pi1951 & ~w8811;
assign w8813 = w8781 & w8785;
assign w8814 = ~w8781 & ~w8785;
assign w8815 = ~w8813 & ~w8814;
assign w8816 = w8793 & w8797;
assign w8817 = ~w8793 & ~w8797;
assign w8818 = ~w8816 & ~w8817;
assign w8819 = pi0346 & ~pi1912;
assign w8820 = ~pi0346 & pi1912;
assign w8821 = ~w8819 & ~w8820;
assign w8822 = pi0411 & ~pi1918;
assign w8823 = ~w8770 & ~w8822;
assign w8824 = w8773 & w8823;
assign w8825 = w2399 & w8821;
assign w8826 = w8824 & w8825;
assign w8827 = w8753 & w8801;
assign w8828 = ~w8821 & w8824;
assign w8829 = ~pi0726 & w8459;
assign w8830 = ~pi1917 & ~pi1921;
assign w8831 = ~pi0780 & w8830;
assign w8832 = ~pi1917 & pi1921;
assign w8833 = ~pi0736 & w8832;
assign w8834 = pi1917 & ~pi1921;
assign w8835 = ~pi0671 & w8834;
assign w8836 = ~w8829 & ~w8831;
assign w8837 = ~w8833 & ~w8835;
assign w8838 = w8836 & w8837;
assign w8839 = ~pi0781 & w8830;
assign w8840 = ~pi0652 & w8832;
assign w8841 = ~pi0727 & w8459;
assign w8842 = ~pi0672 & w8834;
assign w8843 = ~w8839 & ~w8840;
assign w8844 = ~w8841 & ~w8842;
assign w8845 = w8843 & w8844;
assign w8846 = ~pi0783 & w8830;
assign w8847 = ~pi0737 & w8832;
assign w8848 = ~pi0749 & w8834;
assign w8849 = ~pi0639 & w8459;
assign w8850 = ~w8846 & ~w8847;
assign w8851 = ~w8848 & ~w8849;
assign w8852 = w8850 & w8851;
assign w8853 = ~pi0543 & w8832;
assign w8854 = ~pi0530 & w8459;
assign w8855 = ~pi0458 & w8830;
assign w8856 = ~pi0482 & w8834;
assign w8857 = ~w8853 & ~w8854;
assign w8858 = ~w8855 & ~w8856;
assign w8859 = w8857 & w8858;
assign w8860 = ~pi0544 & w8832;
assign w8861 = ~pi0531 & w8459;
assign w8862 = ~pi0483 & w8834;
assign w8863 = ~pi0542 & w8830;
assign w8864 = ~w8860 & ~w8861;
assign w8865 = ~w8862 & ~w8863;
assign w8866 = w8864 & w8865;
assign w8867 = ~pi0729 & w8459;
assign w8868 = ~pi0651 & w8832;
assign w8869 = ~pi0559 & w8834;
assign w8870 = ~pi0637 & w8830;
assign w8871 = ~w8867 & ~w8868;
assign w8872 = ~w8869 & ~w8870;
assign w8873 = w8871 & w8872;
assign w8874 = ~pi0532 & w8459;
assign w8875 = ~pi0484 & w8834;
assign w8876 = ~pi0811 & w8830;
assign w8877 = ~pi0554 & w8832;
assign w8878 = ~w8874 & ~w8875;
assign w8879 = ~w8876 & ~w8877;
assign w8880 = w8878 & w8879;
assign w8881 = ~pi0533 & w8459;
assign w8882 = ~pi0614 & w8830;
assign w8883 = ~pi0485 & w8834;
assign w8884 = ~pi0545 & w8832;
assign w8885 = ~w8881 & ~w8882;
assign w8886 = ~w8883 & ~w8884;
assign w8887 = w8885 & w8886;
assign w8888 = ~pi0534 & w8459;
assign w8889 = ~pi0617 & w8830;
assign w8890 = ~pi0546 & w8832;
assign w8891 = ~pi0486 & w8834;
assign w8892 = ~w8888 & ~w8889;
assign w8893 = ~w8890 & ~w8891;
assign w8894 = w8892 & w8893;
assign w8895 = ~pi0656 & w8830;
assign w8896 = ~pi0535 & w8459;
assign w8897 = ~pi0547 & w8832;
assign w8898 = ~pi0489 & w8834;
assign w8899 = ~w8895 & ~w8896;
assign w8900 = ~w8897 & ~w8898;
assign w8901 = w8899 & w8900;
assign w8902 = w684 & w4921;
assign w8903 = ~pi1993 & ~pi1994;
assign w8904 = w8755 & w8903;
assign w8905 = ~pi1999 & w8827;
assign w8906 = w8904 & w8905;
assign w8907 = ~w8791 & w8798;
assign w8908 = w684 & w7840;
assign w8909 = pi1997 & w8903;
assign w8910 = ~pi1985 & pi1999;
assign w8911 = pi2000 & w8910;
assign w8912 = w8753 & w8909;
assign w8913 = w8911 & w8912;
assign w8914 = w684 & w4939;
assign w8915 = pi1997 & pi1998;
assign w8916 = ~w8904 & w8915;
assign w8917 = ~pi1951 & ~w8916;
assign w8918 = ~pi0734 & w8832;
assign w8919 = ~pi0724 & w8459;
assign w8920 = ~pi0668 & w8834;
assign w8921 = ~pi0641 & w8830;
assign w8922 = ~w8918 & ~w8919;
assign w8923 = ~w8920 & ~w8921;
assign w8924 = w8922 & w8923;
assign w8925 = ~pi0667 & w8834;
assign w8926 = ~pi0660 & w8459;
assign w8927 = ~pi0475 & w8832;
assign w8928 = ~pi0778 & w8830;
assign w8929 = ~w8925 & ~w8926;
assign w8930 = ~w8927 & ~w8928;
assign w8931 = w8929 & w8930;
assign w8932 = ~pi0674 & w8834;
assign w8933 = ~pi0654 & w8832;
assign w8934 = ~pi0779 & w8830;
assign w8935 = ~pi0723 & w8459;
assign w8936 = ~w8932 & ~w8933;
assign w8937 = ~w8934 & ~w8935;
assign w8938 = w8936 & w8937;
assign w8939 = ~pi0735 & w8832;
assign w8940 = ~pi0669 & w8834;
assign w8941 = ~pi0606 & w8830;
assign w8942 = ~pi0725 & w8459;
assign w8943 = ~w8939 & ~w8940;
assign w8944 = ~w8941 & ~w8942;
assign w8945 = w8943 & w8944;
assign w8946 = ~pi0670 & w8834;
assign w8947 = ~pi0605 & w8830;
assign w8948 = ~pi0653 & w8832;
assign w8949 = ~pi0659 & w8459;
assign w8950 = ~w8946 & ~w8947;
assign w8951 = ~w8948 & ~w8949;
assign w8952 = w8950 & w8951;
assign w8953 = ~pi0549 & w8832;
assign w8954 = ~pi0536 & w8459;
assign w8955 = ~pi0624 & w8830;
assign w8956 = ~pi0490 & w8834;
assign w8957 = ~w8953 & ~w8954;
assign w8958 = ~w8955 & ~w8956;
assign w8959 = w8957 & w8958;
assign w8960 = ~pi0492 & w8834;
assign w8961 = ~pi0627 & w8830;
assign w8962 = ~pi0538 & w8459;
assign w8963 = ~pi0551 & w8832;
assign w8964 = ~w8960 & ~w8961;
assign w8965 = ~w8962 & ~w8963;
assign w8966 = w8964 & w8965;
assign w8967 = ~pi0629 & w8830;
assign w8968 = ~pi0552 & w8832;
assign w8969 = ~pi0459 & w8459;
assign w8970 = ~pi0497 & w8834;
assign w8971 = ~w8967 & ~w8968;
assign w8972 = ~w8969 & ~w8970;
assign w8973 = w8971 & w8972;
assign w8974 = ~pi0553 & w8832;
assign w8975 = ~pi0539 & w8459;
assign w8976 = ~pi0632 & w8830;
assign w8977 = ~pi0501 & w8834;
assign w8978 = ~w8974 & ~w8975;
assign w8979 = ~w8976 & ~w8977;
assign w8980 = w8978 & w8979;
assign w8981 = ~pi0744 & w8834;
assign w8982 = ~pi0743 & w8832;
assign w8983 = ~pi0567 & w8459;
assign w8984 = ~pi0603 & w8830;
assign w8985 = ~w8981 & ~w8982;
assign w8986 = ~w8983 & ~w8984;
assign w8987 = w8985 & w8986;
assign w8988 = ~pi0506 & w8834;
assign w8989 = ~pi0555 & w8832;
assign w8990 = ~pi0540 & w8459;
assign w8991 = ~pi0786 & w8830;
assign w8992 = ~w8988 & ~w8989;
assign w8993 = ~w8990 & ~w8991;
assign w8994 = w8992 & w8993;
assign w8995 = ~pi0740 & w8832;
assign w8996 = ~pi0785 & w8830;
assign w8997 = ~pi0562 & w8459;
assign w8998 = ~pi0698 & w8834;
assign w8999 = ~w8995 & ~w8996;
assign w9000 = ~w8997 & ~w8998;
assign w9001 = w8999 & w9000;
assign w9002 = ~pi0753 & w8830;
assign w9003 = ~pi0730 & w8459;
assign w9004 = ~pi0700 & w8834;
assign w9005 = ~pi0741 & w8832;
assign w9006 = ~w9002 & ~w9003;
assign w9007 = ~w9004 & ~w9005;
assign w9008 = w9006 & w9007;
assign w9009 = ~pi0732 & w8459;
assign w9010 = ~pi0787 & w8830;
assign w9011 = ~pi0648 & w8832;
assign w9012 = ~pi0561 & w8834;
assign w9013 = ~w9009 & ~w9010;
assign w9014 = ~w9011 & ~w9012;
assign w9015 = w9013 & w9014;
assign w9016 = ~pi0714 & w8834;
assign w9017 = ~pi0733 & w8459;
assign w9018 = ~pi0788 & w8830;
assign w9019 = ~pi0745 & w8832;
assign w9020 = ~w9016 & ~w9017;
assign w9021 = ~w9018 & ~w9019;
assign w9022 = w9020 & w9021;
assign w9023 = ~pi0655 & w8459;
assign w9024 = ~pi0720 & w8834;
assign w9025 = ~pi0645 & w8832;
assign w9026 = ~pi0752 & w8830;
assign w9027 = ~w9023 & ~w9024;
assign w9028 = ~w9025 & ~w9026;
assign w9029 = w9027 & w9028;
assign w9030 = ~pi0563 & w8834;
assign w9031 = ~pi0568 & w8459;
assign w9032 = ~pi0789 & w8830;
assign w9033 = ~pi0666 & w8832;
assign w9034 = ~w9030 & ~w9031;
assign w9035 = ~w9032 & ~w9033;
assign w9036 = w9034 & w9035;
assign w9037 = ~w8779 & w8786;
assign w9038 = ~pi2000 & w8910;
assign w9039 = pi1993 & w8753;
assign w9040 = w9038 & w9039;
assign w9041 = w8754 & w9040;
assign w9042 = w8623 & w8909;
assign w9043 = w9038 & w9042;
assign w9044 = pi1994 & w8801;
assign w9045 = pi1951 & ~pi1998;
assign w9046 = w9038 & w9045;
assign w9047 = w9044 & w9046;
assign w9048 = w8623 & w8911;
assign w9049 = w9044 & w9048;
assign w9050 = ~pi1994 & ~pi1997;
assign w9051 = w9040 & w9050;
assign w9052 = ~pi1916 & pi1919;
assign w9053 = ~pi0748 & w9052;
assign w9054 = pi1916 & ~pi1919;
assign w9055 = ~pi0692 & w9054;
assign w9056 = ~pi1916 & ~pi1919;
assign w9057 = ~pi0756 & w9056;
assign w9058 = ~pi0707 & w8479;
assign w9059 = ~w9053 & ~w9055;
assign w9060 = ~w9057 & ~w9058;
assign w9061 = w9059 & w9060;
assign w9062 = ~pi0710 & w8479;
assign w9063 = ~pi0758 & w9056;
assign w9064 = ~pi0679 & w9052;
assign w9065 = ~pi0693 & w9054;
assign w9066 = ~w9062 & ~w9063;
assign w9067 = ~w9064 & ~w9065;
assign w9068 = w9066 & w9067;
assign w9069 = ~pi0507 & w9054;
assign w9070 = ~pi0493 & w9052;
assign w9071 = ~pi0519 & w8479;
assign w9072 = ~pi0487 & w9056;
assign w9073 = ~w9069 & ~w9070;
assign w9074 = ~w9071 & ~w9072;
assign w9075 = w9073 & w9074;
assign w9076 = ~pi0520 & w8479;
assign w9077 = ~pi0508 & w9054;
assign w9078 = ~pi0488 & w9056;
assign w9079 = ~pi0494 & w9052;
assign w9080 = ~w9076 & ~w9077;
assign w9081 = ~w9078 & ~w9079;
assign w9082 = w9080 & w9081;
assign w9083 = ~pi0467 & w9054;
assign w9084 = ~pi0521 & w8479;
assign w9085 = ~pi0762 & w9056;
assign w9086 = ~pi0495 & w9052;
assign w9087 = ~w9083 & ~w9084;
assign w9088 = ~w9085 & ~w9086;
assign w9089 = w9087 & w9088;
assign w9090 = ~pi0763 & w9056;
assign w9091 = ~pi0522 & w8479;
assign w9092 = ~pi0510 & w9054;
assign w9093 = ~pi0496 & w9052;
assign w9094 = ~w9090 & ~w9091;
assign w9095 = ~w9092 & ~w9093;
assign w9096 = w9094 & w9095;
assign w9097 = ~pi0764 & w9056;
assign w9098 = ~pi0511 & w9054;
assign w9099 = ~pi0464 & w8479;
assign w9100 = ~pi0470 & w9052;
assign w9101 = ~w9097 & ~w9098;
assign w9102 = ~w9099 & ~w9100;
assign w9103 = w9101 & w9102;
assign w9104 = ~pi0523 & w8479;
assign w9105 = ~pi0512 & w9054;
assign w9106 = ~pi0498 & w9052;
assign w9107 = ~pi0765 & w9056;
assign w9108 = ~w9104 & ~w9105;
assign w9109 = ~w9106 & ~w9107;
assign w9110 = w9108 & w9109;
assign w9111 = ~pi0466 & w9054;
assign w9112 = ~pi0766 & w9056;
assign w9113 = ~pi0524 & w8479;
assign w9114 = ~pi0499 & w9052;
assign w9115 = ~w9111 & ~w9112;
assign w9116 = ~w9113 & ~w9114;
assign w9117 = w9115 & w9116;
assign w9118 = ~pi0469 & w9052;
assign w9119 = ~pi0525 & w8479;
assign w9120 = ~pi0513 & w9054;
assign w9121 = ~pi0767 & w9056;
assign w9122 = ~w9118 & ~w9119;
assign w9123 = ~w9120 & ~w9121;
assign w9124 = w9122 & w9123;
assign w9125 = ~pi0760 & w9056;
assign w9126 = ~pi0680 & w9052;
assign w9127 = ~pi0712 & w8479;
assign w9128 = ~pi0695 & w9054;
assign w9129 = ~w9125 & ~w9126;
assign w9130 = ~w9127 & ~w9128;
assign w9131 = w9129 & w9130;
assign w9132 = ~pi0673 & w8834;
assign w9133 = ~pi0738 & w8832;
assign w9134 = ~pi0728 & w8459;
assign w9135 = ~pi0782 & w8830;
assign w9136 = ~w9132 & ~w9133;
assign w9137 = ~w9134 & ~w9135;
assign w9138 = w9136 & w9137;
assign w9139 = ~pi0514 & w9054;
assign w9140 = ~pi0462 & w8479;
assign w9141 = ~pi0647 & w9056;
assign w9142 = ~pi0500 & w9052;
assign w9143 = ~w9139 & ~w9140;
assign w9144 = ~w9141 & ~w9142;
assign w9145 = w9143 & w9144;
assign w9146 = ~pi0526 & w8479;
assign w9147 = ~pi0502 & w9052;
assign w9148 = ~pi0515 & w9054;
assign w9149 = ~pi0768 & w9056;
assign w9150 = ~w9146 & ~w9147;
assign w9151 = ~w9148 & ~w9149;
assign w9152 = w9150 & w9151;
assign w9153 = ~pi0769 & w9056;
assign w9154 = ~pi0465 & w9054;
assign w9155 = ~pi0468 & w9052;
assign w9156 = ~pi0527 & w8479;
assign w9157 = ~w9153 & ~w9154;
assign w9158 = ~w9155 & ~w9156;
assign w9159 = w9157 & w9158;
assign w9160 = ~pi0770 & w9056;
assign w9161 = ~pi0516 & w9054;
assign w9162 = ~pi0503 & w9052;
assign w9163 = ~pi0528 & w8479;
assign w9164 = ~w9160 & ~w9161;
assign w9165 = ~w9162 & ~w9163;
assign w9166 = w9164 & w9165;
assign w9167 = ~pi0715 & w8479;
assign w9168 = ~pi0683 & w9052;
assign w9169 = ~pi0646 & w9056;
assign w9170 = ~pi0665 & w9054;
assign w9171 = ~w9167 & ~w9168;
assign w9172 = ~w9169 & ~w9170;
assign w9173 = w9171 & w9172;
assign w9174 = ~pi0517 & w9054;
assign w9175 = ~pi0461 & w8479;
assign w9176 = ~pi0504 & w9052;
assign w9177 = ~pi0771 & w9056;
assign w9178 = ~w9174 & ~w9175;
assign w9179 = ~w9176 & ~w9177;
assign w9180 = w9178 & w9179;
assign w9181 = ~pi0529 & w8479;
assign w9182 = ~pi0518 & w9054;
assign w9183 = ~pi0772 & w9056;
assign w9184 = ~pi0505 & w9052;
assign w9185 = ~w9181 & ~w9182;
assign w9186 = ~w9183 & ~w9184;
assign w9187 = w9185 & w9186;
assign w9188 = ~pi0699 & w9054;
assign w9189 = ~pi0684 & w9052;
assign w9190 = ~pi0716 & w8479;
assign w9191 = ~pi0773 & w9056;
assign w9192 = ~w9188 & ~w9189;
assign w9193 = ~w9190 & ~w9191;
assign w9194 = w9192 & w9193;
assign w9195 = ~pi0685 & w9052;
assign w9196 = ~pi0701 & w9054;
assign w9197 = ~pi0642 & w9056;
assign w9198 = ~pi0661 & w8479;
assign w9199 = ~w9195 & ~w9196;
assign w9200 = ~w9197 & ~w9198;
assign w9201 = w9199 & w9200;
assign w9202 = ~pi0774 & w9056;
assign w9203 = ~pi0717 & w8479;
assign w9204 = ~pi0686 & w9052;
assign w9205 = ~pi0664 & w9054;
assign w9206 = ~w9202 & ~w9203;
assign w9207 = ~w9204 & ~w9205;
assign w9208 = w9206 & w9207;
assign w9209 = ~pi0687 & w9052;
assign w9210 = ~pi0775 & w9056;
assign w9211 = ~pi0718 & w8479;
assign w9212 = ~pi0702 & w9054;
assign w9213 = ~w9209 & ~w9210;
assign w9214 = ~w9211 & ~w9212;
assign w9215 = w9213 & w9214;
assign w9216 = ~pi0703 & w9054;
assign w9217 = ~pi0688 & w9052;
assign w9218 = ~pi0776 & w9056;
assign w9219 = ~pi0719 & w8479;
assign w9220 = ~w9216 & ~w9217;
assign w9221 = ~w9218 & ~w9219;
assign w9222 = w9220 & w9221;
assign w9223 = ~pi0689 & w9052;
assign w9224 = ~pi0644 & w9056;
assign w9225 = ~pi0704 & w9054;
assign w9226 = ~pi0722 & w8479;
assign w9227 = ~w9223 & ~w9224;
assign w9228 = ~w9225 & ~w9226;
assign w9229 = w9227 & w9228;
assign w9230 = ~pi0777 & w9056;
assign w9231 = ~pi0739 & w9052;
assign w9232 = ~pi0721 & w8479;
assign w9233 = ~pi0805 & w9054;
assign w9234 = ~w9230 & ~w9231;
assign w9235 = ~w9232 & ~w9233;
assign w9236 = w9234 & w9235;
assign w9237 = ~pi0548 & w8832;
assign w9238 = ~pi0750 & w8830;
assign w9239 = ~pi0471 & w8834;
assign w9240 = ~pi0460 & w8459;
assign w9241 = ~w9237 & ~w9238;
assign w9242 = ~w9239 & ~w9240;
assign w9243 = w9241 & w9242;
assign w9244 = ~pi0537 & w8459;
assign w9245 = ~pi0550 & w8832;
assign w9246 = ~pi0626 & w8830;
assign w9247 = ~pi0491 & w8834;
assign w9248 = ~w9244 & ~w9245;
assign w9249 = ~w9246 & ~w9247;
assign w9250 = w9248 & w9249;
assign w9251 = ~pi0678 & w9052;
assign w9252 = ~pi0709 & w8479;
assign w9253 = ~pi0711 & w9054;
assign w9254 = ~pi0650 & w9056;
assign w9255 = ~w9251 & ~w9252;
assign w9256 = ~w9253 & ~w9254;
assign w9257 = w9255 & w9256;
assign w9258 = ~pi0473 & w8465;
assign w9259 = pi1915 & ~pi1918;
assign w9260 = ~pi0578 & w9259;
assign w9261 = ~pi1915 & ~pi1918;
assign w9262 = ~pi0441 & w9261;
assign w9263 = ~pi1915 & pi1918;
assign w9264 = ~pi0564 & w9263;
assign w9265 = ~w9258 & ~w9260;
assign w9266 = ~w9262 & ~w9264;
assign w9267 = w9265 & w9266;
assign w9268 = ~pi0442 & w9261;
assign w9269 = ~pi0565 & w9263;
assign w9270 = ~pi0596 & w8465;
assign w9271 = ~pi0579 & w9259;
assign w9272 = ~w9268 & ~w9269;
assign w9273 = ~w9270 & ~w9271;
assign w9274 = w9272 & w9273;
assign w9275 = ~pi0593 & w8465;
assign w9276 = ~pi0443 & w9261;
assign w9277 = ~pi0566 & w9263;
assign w9278 = ~pi0580 & w9259;
assign w9279 = ~w9275 & ~w9276;
assign w9280 = ~w9277 & ~w9278;
assign w9281 = w9279 & w9280;
assign w9282 = ~pi0444 & w9261;
assign w9283 = ~pi0400 & w9263;
assign w9284 = ~pi0586 & w9259;
assign w9285 = ~pi0594 & w8465;
assign w9286 = ~w9282 & ~w9283;
assign w9287 = ~w9284 & ~w9285;
assign w9288 = w9286 & w9287;
assign w9289 = ~pi0581 & w9259;
assign w9290 = ~pi0445 & w9261;
assign w9291 = ~pi0401 & w9263;
assign w9292 = ~pi0474 & w8465;
assign w9293 = ~w9289 & ~w9290;
assign w9294 = ~w9291 & ~w9292;
assign w9295 = w9293 & w9294;
assign w9296 = ~pi0784 & w8830;
assign w9297 = ~pi0556 & w8832;
assign w9298 = ~pi0509 & w8834;
assign w9299 = ~pi0541 & w8459;
assign w9300 = ~w9296 & ~w9297;
assign w9301 = ~w9298 & ~w9299;
assign w9302 = w9300 & w9301;
assign w9303 = ~pi0582 & w9259;
assign w9304 = ~pi0569 & w9263;
assign w9305 = ~pi0472 & w8465;
assign w9306 = ~pi0446 & w9261;
assign w9307 = ~w9303 & ~w9304;
assign w9308 = ~w9305 & ~w9306;
assign w9309 = w9307 & w9308;
assign w9310 = ~pi0447 & w9261;
assign w9311 = ~pi0595 & w8465;
assign w9312 = ~pi0476 & w9263;
assign w9313 = ~pi0583 & w9259;
assign w9314 = ~w9310 & ~w9311;
assign w9315 = ~w9312 & ~w9313;
assign w9316 = w9314 & w9315;
assign w9317 = ~pi0402 & w9263;
assign w9318 = ~pi0607 & w9261;
assign w9319 = ~pi0584 & w9259;
assign w9320 = ~pi0407 & w8465;
assign w9321 = ~w9317 & ~w9318;
assign w9322 = ~w9319 & ~w9320;
assign w9323 = w9321 & w9322;
assign w9324 = ~pi0638 & w9261;
assign w9325 = ~pi0585 & w9263;
assign w9326 = ~pi0403 & w9259;
assign w9327 = ~pi0408 & w8465;
assign w9328 = ~w9324 & ~w9325;
assign w9329 = ~w9326 & ~w9327;
assign w9330 = w9328 & w9329;
assign w9331 = ~pi0371 & w9259;
assign w9332 = ~pi0385 & w8465;
assign w9333 = ~pi0357 & w9263;
assign w9334 = ~pi0355 & w9261;
assign w9335 = ~w9331 & ~w9332;
assign w9336 = ~w9333 & ~w9334;
assign w9337 = w9335 & w9336;
assign w9338 = ~pi0386 & w8465;
assign w9339 = ~pi0358 & w9263;
assign w9340 = ~pi0372 & w9259;
assign w9341 = ~pi0356 & w9261;
assign w9342 = ~w9338 & ~w9339;
assign w9343 = ~w9340 & ~w9341;
assign w9344 = w9342 & w9343;
assign w9345 = ~pi0560 & w8834;
assign w9346 = ~pi0634 & w8830;
assign w9347 = ~pi0742 & w8832;
assign w9348 = ~pi0731 & w8459;
assign w9349 = ~w9345 & ~w9346;
assign w9350 = ~w9347 & ~w9348;
assign w9351 = w9349 & w9350;
assign w9352 = ~pi0570 & w9263;
assign w9353 = ~pi0404 & w9259;
assign w9354 = ~pi0448 & w9261;
assign w9355 = ~pi0600 & w8465;
assign w9356 = ~w9352 & ~w9353;
assign w9357 = ~w9354 & ~w9355;
assign w9358 = w9356 & w9357;
assign w9359 = ~pi0373 & w9259;
assign w9360 = ~pi0608 & w9261;
assign w9361 = ~pi0387 & w8465;
assign w9362 = ~pi0359 & w9263;
assign w9363 = ~w9359 & ~w9360;
assign w9364 = ~w9361 & ~w9362;
assign w9365 = w9363 & w9364;
assign w9366 = ~pi0388 & w8465;
assign w9367 = ~pi0360 & w9263;
assign w9368 = ~pi0374 & w9259;
assign w9369 = ~pi0609 & w9261;
assign w9370 = ~w9366 & ~w9367;
assign w9371 = ~w9368 & ~w9369;
assign w9372 = w9370 & w9371;
assign w9373 = ~pi0361 & w9263;
assign w9374 = ~pi0610 & w9261;
assign w9375 = ~pi0375 & w9259;
assign w9376 = ~pi0389 & w8465;
assign w9377 = ~w9373 & ~w9374;
assign w9378 = ~w9375 & ~w9376;
assign w9379 = w9377 & w9378;
assign w9380 = ~pi0362 & w9263;
assign w9381 = ~pi0390 & w8465;
assign w9382 = ~pi0611 & w9261;
assign w9383 = ~pi0376 & w9259;
assign w9384 = ~w9380 & ~w9381;
assign w9385 = ~w9382 & ~w9383;
assign w9386 = w9384 & w9385;
assign w9387 = ~pi0363 & w9263;
assign w9388 = ~pi0377 & w9259;
assign w9389 = ~pi0391 & w8465;
assign w9390 = ~pi0612 & w9261;
assign w9391 = ~w9387 & ~w9388;
assign w9392 = ~w9389 & ~w9390;
assign w9393 = w9391 & w9392;
assign w9394 = ~pi0613 & w9261;
assign w9395 = ~pi0378 & w9259;
assign w9396 = ~pi0364 & w9263;
assign w9397 = ~pi0392 & w8465;
assign w9398 = ~w9394 & ~w9395;
assign w9399 = ~w9396 & ~w9397;
assign w9400 = w9398 & w9399;
assign w9401 = ~pi0615 & w9261;
assign w9402 = ~pi0379 & w9259;
assign w9403 = ~pi0365 & w9263;
assign w9404 = ~pi0393 & w8465;
assign w9405 = ~w9401 & ~w9402;
assign w9406 = ~w9403 & ~w9404;
assign w9407 = w9405 & w9406;
assign w9408 = ~pi0380 & w9259;
assign w9409 = ~pi0366 & w9263;
assign w9410 = ~pi0616 & w9261;
assign w9411 = ~pi0394 & w8465;
assign w9412 = ~w9408 & ~w9409;
assign w9413 = ~w9410 & ~w9411;
assign w9414 = w9412 & w9413;
assign w9415 = ~pi0618 & w9261;
assign w9416 = ~pi0395 & w8465;
assign w9417 = ~pi0367 & w9263;
assign w9418 = ~pi0381 & w9259;
assign w9419 = ~w9415 & ~w9416;
assign w9420 = ~w9417 & ~w9418;
assign w9421 = w9419 & w9420;
assign w9422 = ~pi0382 & w9259;
assign w9423 = ~pi0619 & w9261;
assign w9424 = ~pi0396 & w8465;
assign w9425 = ~pi0368 & w9263;
assign w9426 = ~w9422 & ~w9423;
assign w9427 = ~w9424 & ~w9425;
assign w9428 = w9426 & w9427;
assign w9429 = ~pi0571 & w9263;
assign w9430 = ~pi0597 & w8465;
assign w9431 = ~pi0587 & w9259;
assign w9432 = ~pi0620 & w9261;
assign w9433 = ~w9429 & ~w9430;
assign w9434 = ~w9431 & ~w9432;
assign w9435 = w9433 & w9434;
assign w9436 = ~pi0369 & w9263;
assign w9437 = ~pi0383 & w9259;
assign w9438 = ~pi0621 & w9261;
assign w9439 = ~pi0397 & w8465;
assign w9440 = ~w9436 & ~w9437;
assign w9441 = ~w9438 & ~w9439;
assign w9442 = w9440 & w9441;
assign w9443 = ~pi0370 & w9263;
assign w9444 = ~pi0398 & w8465;
assign w9445 = ~pi0622 & w9261;
assign w9446 = ~pi0384 & w9259;
assign w9447 = ~w9443 & ~w9444;
assign w9448 = ~w9445 & ~w9446;
assign w9449 = w9447 & w9448;
assign w9450 = ~pi0572 & w9263;
assign w9451 = ~pi0598 & w8465;
assign w9452 = ~pi0588 & w9259;
assign w9453 = ~pi0623 & w9261;
assign w9454 = ~w9450 & ~w9451;
assign w9455 = ~w9452 & ~w9453;
assign w9456 = w9454 & w9455;
assign w9457 = ~pi0590 & w9259;
assign w9458 = ~pi0625 & w9261;
assign w9459 = ~pi0599 & w8465;
assign w9460 = ~pi0573 & w9263;
assign w9461 = ~w9457 & ~w9458;
assign w9462 = ~w9459 & ~w9460;
assign w9463 = w9461 & w9462;
assign w9464 = ~pi0409 & w8465;
assign w9465 = ~pi0574 & w9263;
assign w9466 = ~pi0591 & w9259;
assign w9467 = ~pi0604 & w9261;
assign w9468 = ~w9464 & ~w9465;
assign w9469 = ~w9466 & ~w9467;
assign w9470 = w9468 & w9469;
assign w9471 = ~pi0589 & w9259;
assign w9472 = ~pi0628 & w9261;
assign w9473 = ~pi0410 & w8465;
assign w9474 = ~pi0477 & w9263;
assign w9475 = ~w9471 & ~w9472;
assign w9476 = ~w9473 & ~w9474;
assign w9477 = w9475 & w9476;
assign w9478 = ~pi0405 & w9259;
assign w9479 = ~pi0630 & w9261;
assign w9480 = ~pi0575 & w9263;
assign w9481 = ~pi0399 & w8465;
assign w9482 = ~w9478 & ~w9479;
assign w9483 = ~w9480 & ~w9481;
assign w9484 = w9482 & w9483;
assign w9485 = ~pi0557 & w8465;
assign w9486 = ~pi0631 & w9261;
assign w9487 = ~pi0576 & w9263;
assign w9488 = ~pi0406 & w9259;
assign w9489 = ~w9485 & ~w9486;
assign w9490 = ~w9487 & ~w9488;
assign w9491 = w9489 & w9490;
assign w9492 = ~pi0577 & w9263;
assign w9493 = ~pi0633 & w9261;
assign w9494 = ~pi0592 & w9259;
assign w9495 = ~pi0558 & w8465;
assign w9496 = ~w9492 & ~w9493;
assign w9497 = ~w9494 & ~w9495;
assign w9498 = w9496 & w9497;
assign w9499 = ~pi0747 & w9052;
assign w9500 = ~pi0759 & w9056;
assign w9501 = ~pi0663 & w8479;
assign w9502 = ~pi0694 & w9054;
assign w9503 = ~w9499 & ~w9500;
assign w9504 = ~w9501 & ~w9502;
assign w9505 = w9503 & w9504;
assign w9506 = ~pi0713 & w8479;
assign w9507 = ~pi0696 & w9054;
assign w9508 = ~pi0649 & w9056;
assign w9509 = ~pi0681 & w9052;
assign w9510 = ~w9506 & ~w9507;
assign w9511 = ~w9508 & ~w9509;
assign w9512 = w9510 & w9511;
assign w9513 = ~pi0690 & w9054;
assign w9514 = ~pi0675 & w9052;
assign w9515 = ~pi0754 & w9056;
assign w9516 = ~pi0705 & w8479;
assign w9517 = ~w9513 & ~w9514;
assign w9518 = ~w9515 & ~w9516;
assign w9519 = w9517 & w9518;
assign w9520 = ~pi0757 & w9056;
assign w9521 = ~pi0708 & w8479;
assign w9522 = ~pi0677 & w9052;
assign w9523 = ~pi0658 & w9054;
assign w9524 = ~w9520 & ~w9521;
assign w9525 = ~w9522 & ~w9523;
assign w9526 = w9524 & w9525;
assign w9527 = ~pi0691 & w9054;
assign w9528 = ~pi0676 & w9052;
assign w9529 = ~pi0706 & w8479;
assign w9530 = ~pi0755 & w9056;
assign w9531 = ~w9527 & ~w9528;
assign w9532 = ~w9529 & ~w9530;
assign w9533 = w9531 & w9532;
assign w9534 = ~pi0662 & w8479;
assign w9535 = ~pi0697 & w9054;
assign w9536 = ~pi0761 & w9056;
assign w9537 = ~pi0682 & w9052;
assign w9538 = ~w9534 & ~w9535;
assign w9539 = ~w9536 & ~w9537;
assign w9540 = w9538 & w9539;
assign w9541 = w683 & w8806;
assign w9542 = pi2163 & ~pi2180;
assign w9543 = ~pi2163 & pi2180;
assign w9544 = ~w9542 & ~w9543;
assign w9545 = pi0873 & pi0878;
assign w9546 = ~pi0873 & pi2143;
assign w9547 = ~w9545 & ~w9546;
assign w9548 = pi0478 & pi0873;
assign w9549 = ~pi0873 & pi2144;
assign w9550 = ~w9548 & ~w9549;
assign w9551 = pi0210 & pi0873;
assign w9552 = ~pi0873 & pi2145;
assign w9553 = ~w9551 & ~w9552;
assign w9554 = pi0873 & pi1923;
assign w9555 = ~pi0873 & pi2146;
assign w9556 = ~w9554 & ~w9555;
assign w9557 = pi0869 & pi0873;
assign w9558 = ~pi0873 & pi2147;
assign w9559 = ~w9557 & ~w9558;
assign w9560 = pi0194 & pi0873;
assign w9561 = ~pi0873 & pi2148;
assign w9562 = ~w9560 & ~w9561;
assign w9563 = pi0336 & pi0873;
assign w9564 = ~pi0873 & pi2149;
assign w9565 = ~w9563 & ~w9564;
assign w9566 = pi0190 & pi0873;
assign w9567 = ~pi0873 & pi2150;
assign w9568 = ~w9566 & ~w9567;
assign w9569 = pi0873 & pi0948;
assign w9570 = ~pi0873 & pi2151;
assign w9571 = ~w9569 & ~w9570;
assign w9572 = pi0817 & pi0873;
assign w9573 = ~pi0873 & pi2152;
assign w9574 = ~w9572 & ~w9573;
assign w9575 = pi0234 & pi0873;
assign w9576 = ~pi0873 & pi2153;
assign w9577 = ~w9575 & ~w9576;
assign w9578 = pi0205 & pi0873;
assign w9579 = ~pi0873 & pi2154;
assign w9580 = ~w9578 & ~w9579;
assign w9581 = pi0873 & pi1885;
assign w9582 = ~pi0873 & pi2155;
assign w9583 = ~w9581 & ~w9582;
assign w9584 = pi0873 & pi1932;
assign w9585 = ~pi0873 & pi2156;
assign w9586 = ~w9584 & ~w9585;
assign w9587 = pi0873 & pi0906;
assign w9588 = ~pi0873 & pi2157;
assign w9589 = ~w9587 & ~w9588;
assign w9590 = ~w5018 & ~w5019;
assign w9591 = pi0873 & pi1851;
assign w9592 = ~pi0873 & pi2160;
assign w9593 = ~w9591 & ~w9592;
assign w9594 = pi1035 & pi1168;
assign w9595 = w9594 & pi0329;
assign w9596 = ~w9595 & ~pi0198;
assign w9597 = pi1176 & pi1181;
assign w9598 = w9597 & pi0330;
assign w9599 = ~w9598 & ~pi0199;
assign w9600 = pi1164 & pi1185;
assign w9601 = w9600 & pi0341;
assign w9602 = ~w9601 & ~pi0201;
assign w9603 = pi1169 & pi1762;
assign w9604 = w9603 & pi0342;
assign w9605 = ~w9604 & ~pi0202;
assign w9606 = pi1839 & pi1848;
assign w9607 = w9606 & pi0343;
assign w9608 = ~w9607 & ~pi0203;
assign w9609 = pi1838 & pi1843;
assign w9610 = w9609 & pi0344;
assign w9611 = ~w9610 & ~pi0204;
assign w9612 = pi1035 & pi0214;
assign w9613 = pi1035 & ~w2284;
assign w9614 = pi1169 & w610;
assign w9615 = ~pi0238 & pi1169;
assign w9616 = ~w9614 & ~pi0215;
assign w9617 = pi1838 & pi0216;
assign w9618 = pi1838 & ~w865;
assign w9619 = pi1164 & pi0217;
assign w9620 = pi1164 & ~w819;
assign w9621 = pi1176 & pi0218;
assign w9622 = pi1176 & ~w721;
assign w9623 = pi1839 & pi0219;
assign w9624 = pi1839 & ~w771;
assign w9625 = ~w863 & ~pi0220;
assign w9626 = w863 & pi0220;
assign w9627 = pi1838 & pi0220;
assign w9628 = pi1838 & ~w9625;
assign w9629 = ~w813 & ~pi0221;
assign w9630 = w813 & pi0221;
assign w9631 = pi1164 & pi0221;
assign w9632 = pi1164 & ~w9629;
assign w9633 = ~w725 & ~pi0222;
assign w9634 = w725 & pi0222;
assign w9635 = pi1176 & pi0222;
assign w9636 = pi1176 & ~w9633;
assign w9637 = ~w773 & ~pi0223;
assign w9638 = w773 & pi0223;
assign w9639 = pi1839 & pi0223;
assign w9640 = pi1839 & ~w9637;
assign w9641 = ~pi0224 & pi1838;
assign w9642 = ~pi0225 & pi1164;
assign w9643 = ~pi0226 & pi1839;
assign w9644 = ~pi0227 & pi1176;
assign w9645 = ~pi0236 & pi1035;
assign w9646 = ~w2282 & ~pi0237;
assign w9647 = w2282 & pi0237;
assign w9648 = pi1035 & pi0237;
assign w9649 = pi1035 & ~w9646;
assign w9650 = pi1169 & w715;
assign w9651 = ~pi1078 & pi1176;
assign w9652 = pi1078 & pi1176;
assign w9653 = ~w720 & ~w733;
assign w9654 = ~w720 & ~w753;
assign w9655 = ~pi1079 & pi1839;
assign w9656 = pi1079 & pi1839;
assign w9657 = ~w766 & ~w779;
assign w9658 = ~w766 & ~w799;
assign w9659 = ~pi1075 & pi1164;
assign w9660 = pi1075 & pi1164;
assign w9661 = ~w812 & ~w825;
assign w9662 = ~w827 & ~w845;
assign w9663 = ~pi1080 & pi1838;
assign w9664 = pi1080 & pi1838;
assign w9665 = ~w858 & ~w871;
assign w9666 = ~w858 & ~w891;
assign w9667 = ~w623 & w935;
assign w9668 = ~w631 & w939;
assign w9669 = ~w639 & ~pi0262;
assign w9670 = w639 & pi0262;
assign w9671 = ~w647 & ~pi0263;
assign w9672 = w647 & pi0263;
assign w9673 = ~w735 & ~w959;
assign w9674 = ~w967 & ~w996;
assign w9675 = ~w967 & ~w1032;
assign w9676 = ~w967 & ~w1054;
assign w9677 = ~w720 & ~w1076;
assign w9678 = ~w967 & ~w1098;
assign w9679 = ~w735 & ~w1120;
assign w9680 = ~w735 & ~w1149;
assign w9681 = ~w720 & ~w1178;
assign w9682 = ~w735 & ~w1193;
assign w9683 = ~w735 & ~w1207;
assign w9684 = ~w720 & ~w1215;
assign w9685 = ~w967 & ~w1232;
assign w9686 = ~w967 & ~w1240;
assign w9687 = ~w720 & ~w1254;
assign w9688 = ~w967 & ~w1269;
assign w9689 = ~w1286 & ~w1285;
assign w9690 = ~w766 & ~w1322;
assign w9691 = ~w781 & ~w1358;
assign w9692 = ~w1286 & ~w1380;
assign w9693 = ~w766 & ~w1402;
assign w9694 = ~w766 & ~w1424;
assign w9695 = ~w1286 & ~w1453;
assign w9696 = ~w781 & ~w1468;
assign w9697 = ~w766 & ~w1490;
assign w9698 = ~w781 & ~w1512;
assign w9699 = ~w1286 & ~w1526;
assign w9700 = ~w1286 & ~w1541;
assign w9701 = ~w766 & ~w1558;
assign w9702 = ~w781 & ~w1566;
assign w9703 = ~w766 & ~w1580;
assign w9704 = ~w766 & ~w1595;
assign w9705 = w631 & w939;
assign w9706 = ~w827 & ~w1609;
assign w9707 = ~w827 & ~w1646;
assign w9708 = ~w812 & ~w1675;
assign w9709 = ~w827 & ~w1704;
assign w9710 = ~w812 & ~w1726;
assign w9711 = ~w812 & ~w1748;
assign w9712 = ~w812 & ~w1770;
assign w9713 = ~w827 & ~w1799;
assign w9714 = w623 & w935;
assign w9715 = ~w934 & ~w1821;
assign w9716 = ~w827 & ~w1858;
assign w9717 = ~w873 & ~w1880;
assign w9718 = ~w934 & ~w1909;
assign w9719 = ~w827 & ~w1931;
assign w9720 = ~w873 & ~w1946;
assign w9721 = ~w858 & ~w1975;
assign w9722 = ~w1626 & ~w1990;
assign w9723 = ~w858 & ~w2012;
assign w9724 = ~w812 & ~w2027;
assign w9725 = ~w858 & ~w2042;
assign w9726 = ~w812 & ~w2071;
assign w9727 = ~w858 & ~w2086;
assign w9728 = ~w827 & ~w2101;
assign w9729 = ~w858 & ~w2116;
assign w9730 = ~w1626 & ~w2131;
assign w9731 = ~w858 & ~w2146;
assign w9732 = ~w812 & ~w2161;
assign w9733 = ~w858 & ~w2183;
assign w9734 = ~w858 & ~w2198;
assign w9735 = ~w934 & ~w2206;
assign w9736 = ~w934 & ~w2214;
assign w9737 = ~w873 & ~w2222;
assign w9738 = ~w858 & ~w2237;
assign w9739 = pi1150 & pi1128;
assign w9740 = w9739 & pi0865;
assign w9741 = ~w9740 & ~pi0332;
assign w9742 = ~pi1076 & pi1035;
assign w9743 = pi1076 & pi1035;
assign w9744 = ~w2281 & ~w2294;
assign w9745 = ~pi1077 & pi1169;
assign w9746 = pi1077 & pi1169;
assign w9747 = ~w2309 & ~w2320;
assign w9748 = ~w2309 & ~w2340;
assign w9749 = ~w2281 & ~w2358;
assign w9750 = w604 & w2383;
assign w9751 = ~w2373 & ~w2374;
assign w9752 = pi0411 & pi0412;
assign w9753 = ~w9752 & ~pi0346;
assign w9754 = w9752 & pi0346;
assign w9755 = pi1150 & pi0346;
assign w9756 = pi1150 & ~w9753;
assign w9757 = pi1145 & pi1161;
assign w9758 = w9757 & pi0874;
assign w9759 = ~w9758 & ~pi0347;
assign w9760 = pi1036 & pi1149;
assign w9761 = w9760 & pi0875;
assign w9762 = ~w9761 & ~pi0348;
assign w9763 = ~w604 & w2383;
assign w9764 = ~w611 & w2442;
assign w9765 = ~pi0411 & ~pi0412;
assign w9766 = ~w9765 & ~pi0355;
assign w9767 = ~w9765 & ~pi0356;
assign w9768 = pi0411 & ~pi0412;
assign w9769 = ~w9768 & ~pi0357;
assign w9770 = ~w9768 & ~pi0358;
assign w9771 = w9768 & w2398;
assign w9772 = w9771 & pi0947;
assign w9773 = ~w9768 & ~pi0359;
assign w9774 = w9771 & pi0923;
assign w9775 = ~w9768 & ~pi0360;
assign w9776 = w9771 & pi0877;
assign w9777 = ~w9768 & ~pi0361;
assign w9778 = w9771 & pi0871;
assign w9779 = ~w9768 & ~pi0362;
assign w9780 = w9771 & pi0814;
assign w9781 = ~w9768 & ~pi0363;
assign w9782 = w9771 & pi0480;
assign w9783 = ~w9768 & ~pi0364;
assign w9784 = w9771 & pi0335;
assign w9785 = ~w9768 & ~pi0365;
assign w9786 = w9771 & pi0233;
assign w9787 = ~w9768 & ~pi0366;
assign w9788 = w9771 & pi0213;
assign w9789 = ~w9768 & ~pi0367;
assign w9790 = w9771 & pi0208;
assign w9791 = ~w9768 & ~pi0368;
assign w9792 = w9771 & pi0197;
assign w9793 = ~w9768 & ~pi0369;
assign w9794 = w9771 & pi0193;
assign w9795 = ~pi0411 & pi0412;
assign w9796 = ~w9795 & ~pi0371;
assign w9797 = ~w9795 & ~pi0372;
assign w9798 = w9795 & w2398;
assign w9799 = w9798 & pi0947;
assign w9800 = ~w9795 & ~pi0373;
assign w9801 = w9798 & pi0923;
assign w9802 = ~w9795 & ~pi0374;
assign w9803 = w9798 & pi0877;
assign w9804 = ~w9795 & ~pi0375;
assign w9805 = w9798 & pi0871;
assign w9806 = ~w9795 & ~pi0376;
assign w9807 = w9798 & pi0814;
assign w9808 = ~w9795 & ~pi0377;
assign w9809 = w9798 & pi0480;
assign w9810 = ~w9795 & ~pi0378;
assign w9811 = w9798 & pi0335;
assign w9812 = ~w9795 & ~pi0379;
assign w9813 = w9798 & pi0233;
assign w9814 = ~w9795 & ~pi0380;
assign w9815 = w9798 & pi0213;
assign w9816 = ~w9795 & ~pi0381;
assign w9817 = w9798 & pi0208;
assign w9818 = ~w9795 & ~pi0382;
assign w9819 = w9798 & pi0197;
assign w9820 = ~w9795 & ~pi0383;
assign w9821 = w9798 & pi0193;
assign w9822 = ~w9752 & ~pi0385;
assign w9823 = ~w9752 & ~pi0386;
assign w9824 = w9752 & w2398;
assign w9825 = w9824 & pi0947;
assign w9826 = ~w9752 & ~pi0387;
assign w9827 = w9824 & pi0923;
assign w9828 = ~w9752 & ~pi0388;
assign w9829 = w9824 & pi0877;
assign w9830 = ~w9752 & ~pi0389;
assign w9831 = w9824 & pi0871;
assign w9832 = ~w9752 & ~pi0390;
assign w9833 = w9824 & pi0814;
assign w9834 = ~w9752 & ~pi0391;
assign w9835 = w9824 & pi0480;
assign w9836 = ~w9752 & ~pi0392;
assign w9837 = w9824 & pi0335;
assign w9838 = ~w9752 & ~pi0393;
assign w9839 = w9824 & pi0233;
assign w9840 = ~w9752 & ~pi0394;
assign w9841 = w9824 & pi0213;
assign w9842 = ~w9752 & ~pi0395;
assign w9843 = w9824 & pi0208;
assign w9844 = ~w9752 & ~pi0396;
assign w9845 = w9824 & pi0197;
assign w9846 = ~w9752 & ~pi0397;
assign w9847 = w9824 & pi0193;
assign w9848 = ~w9752 & ~pi0399;
assign w9849 = ~w9768 & ~pi0400;
assign w9850 = ~w9768 & ~pi0401;
assign w9851 = ~w9768 & ~pi0402;
assign w9852 = ~w9795 & ~pi0403;
assign w9853 = ~w9795 & ~pi0404;
assign w9854 = ~w9795 & ~pi0405;
assign w9855 = ~w9795 & ~pi0406;
assign w9856 = ~w9752 & ~pi0407;
assign w9857 = ~w9752 & ~pi0408;
assign w9858 = ~w9752 & ~pi0409;
assign w9859 = ~w9752 & ~pi0410;
assign w9860 = ~pi0411 & pi1150;
assign w9861 = ~w2296 & ~w2682;
assign w9862 = ~w2281 & ~w2718;
assign w9863 = ~w2296 & ~w2754;
assign w9864 = ~w2296 & ~w2783;
assign w9865 = ~w2281 & ~w2798;
assign w9866 = ~w2296 & ~w2813;
assign w9867 = ~w2296 & ~w2842;
assign w9868 = ~w2296 & ~w2857;
assign w9869 = ~w2296 & ~w2879;
assign w9870 = ~w2281 & ~w2901;
assign w9871 = ~w2384 & ~w2916;
assign w9872 = ~w2281 & ~w2931;
assign w9873 = ~w2281 & ~w2939;
assign w9874 = ~w2281 & ~w2947;
assign w9875 = ~w2281 & ~w2962;
assign w9876 = w611 & w2442;
assign w9877 = ~w2441 & ~w2984;
assign w9878 = ~w2309 & ~w3021;
assign w9879 = ~w2441 & ~w3050;
assign w9880 = ~w2322 & ~w3079;
assign w9881 = ~w2441 & ~w3094;
assign w9882 = ~w2322 & ~w3130;
assign w9883 = ~w2322 & ~w3152;
assign w9884 = ~w2322 & ~w3174;
assign w9885 = ~w2322 & ~w3203;
assign w9886 = ~w3001 & ~w3211;
assign w9887 = ~w2441 & ~w3226;
assign w9888 = ~w2309 & ~w3234;
assign w9889 = ~w2322 & ~w3249;
assign w9890 = ~w9765 & ~pi0441;
assign w9891 = ~w9765 & ~pi0442;
assign w9892 = ~w9765 & ~pi0443;
assign w9893 = ~w9765 & ~pi0444;
assign w9894 = ~w9765 & ~pi0445;
assign w9895 = ~w9765 & ~pi0446;
assign w9896 = ~w9765 & ~pi0447;
assign w9897 = ~w9765 & ~pi0448;
assign w9898 = ~pi0836 & pi0449;
assign w9899 = ~pi1075 & ~pi1907;
assign w9900 = ~pi1078 & ~pi1904;
assign w9901 = ~pi1079 & ~pi1909;
assign w9902 = ~pi1080 & ~pi1910;
assign w9903 = ~w2322 & ~w3325;
assign w9904 = ~w2441 & ~w3333;
assign w9905 = ~w2309 & ~w3348;
assign w9906 = ~pi0601 & ~pi0602;
assign w9907 = ~w9906 & ~pi0458;
assign w9908 = pi0601 & pi0602;
assign w9909 = w9908 & w3363;
assign w9910 = w9909 & pi0212;
assign w9911 = ~w9908 & ~pi0459;
assign w9912 = w9909 & pi0819;
assign w9913 = ~w9908 & ~pi0460;
assign w9914 = pi0843 & pi0746;
assign w9915 = w9914 & w3383;
assign w9916 = w9915 & pi0195;
assign w9917 = ~w9914 & ~pi0461;
assign w9918 = w9915 & pi0333;
assign w9919 = ~w9914 & ~pi0462;
assign w9920 = ~w9908 & ~pi0463;
assign w9921 = w9908 & pi0463;
assign w9922 = pi1036 & pi0463;
assign w9923 = pi1036 & ~w9920;
assign w9924 = w9915 & pi0883;
assign w9925 = ~w9914 & ~pi0464;
assign w9926 = ~pi0843 & pi0746;
assign w9927 = w9926 & w3383;
assign w9928 = w9927 & pi0211;
assign w9929 = ~w9926 & ~pi0465;
assign w9930 = w9927 & pi0818;
assign w9931 = ~w9926 & ~pi0466;
assign w9932 = w9927 & pi0951;
assign w9933 = ~w9926 & ~pi0467;
assign w9934 = pi0843 & ~pi0746;
assign w9935 = w9934 & w3383;
assign w9936 = w9935 & pi0211;
assign w9937 = ~w9934 & ~pi0468;
assign w9938 = w9935 & pi0481;
assign w9939 = ~w9934 & ~pi0469;
assign w9940 = w9935 & pi0883;
assign w9941 = ~w9934 & ~pi0470;
assign w9942 = ~pi0601 & pi0602;
assign w9943 = w3363 & pi0819;
assign w9944 = ~w9942 & ~pi0471;
assign w9945 = ~w9752 & ~pi0472;
assign w9946 = ~w9752 & ~pi0473;
assign w9947 = ~w9752 & ~pi0474;
assign w9948 = pi0601 & ~pi0602;
assign w9949 = ~w9948 & ~pi0475;
assign w9950 = ~w9768 & ~pi0476;
assign w9951 = ~w9768 & ~pi0477;
assign w9952 = ~w9942 & ~pi0482;
assign w9953 = ~w9942 & ~pi0483;
assign w9954 = w3363 & pi0950;
assign w9955 = ~w9942 & ~pi0484;
assign w9956 = w3363 & pi0915;
assign w9957 = ~w9942 & ~pi0485;
assign w9958 = w3363 & pi0882;
assign w9959 = ~w9942 & ~pi0486;
assign w9960 = ~pi0843 & ~pi0746;
assign w9961 = ~w9960 & ~pi0487;
assign w9962 = ~w9960 & ~pi0488;
assign w9963 = w3363 & pi0866;
assign w9964 = ~w9942 & ~pi0489;
assign w9965 = w3363 & pi0479;
assign w9966 = ~w9942 & ~pi0490;
assign w9967 = w3363 & pi0334;
assign w9968 = ~w9942 & ~pi0491;
assign w9969 = w3363 & pi0235;
assign w9970 = ~w9942 & ~pi0492;
assign w9971 = ~w9934 & ~pi0493;
assign w9972 = ~w9934 & ~pi0494;
assign w9973 = w9935 & pi0951;
assign w9974 = ~w9934 & ~pi0495;
assign w9975 = w9935 & pi0916;
assign w9976 = ~w9934 & ~pi0496;
assign w9977 = w3363 & pi0212;
assign w9978 = ~w9942 & ~pi0497;
assign w9979 = w9935 & pi0870;
assign w9980 = ~w9934 & ~pi0498;
assign w9981 = w9935 & pi0818;
assign w9982 = ~w9934 & ~pi0499;
assign w9983 = w9935 & pi0333;
assign w9984 = ~w9934 & ~pi0500;
assign w9985 = w3363 & pi0207;
assign w9986 = ~w9942 & ~pi0501;
assign w9987 = w9935 & pi0231;
assign w9988 = ~w9934 & ~pi0502;
assign w9989 = w9935 & pi0206;
assign w9990 = ~w9934 & ~pi0503;
assign w9991 = w9935 & pi0195;
assign w9992 = ~w9934 & ~pi0504;
assign w9993 = w9935 & pi0191;
assign w9994 = w3363 & pi0196;
assign w9995 = ~w9942 & ~pi0506;
assign w9996 = ~w9926 & ~pi0507;
assign w9997 = ~w9926 & ~pi0508;
assign w9998 = w3363 & pi0192;
assign w9999 = w9927 & pi0916;
assign w10000 = ~w9926 & ~pi0510;
assign w10001 = w9927 & pi0883;
assign w10002 = ~w9926 & ~pi0511;
assign w10003 = w9927 & pi0870;
assign w10004 = ~w9926 & ~pi0512;
assign w10005 = w9927 & pi0481;
assign w10006 = ~w9926 & ~pi0513;
assign w10007 = w9927 & pi0333;
assign w10008 = ~w9926 & ~pi0514;
assign w10009 = w9927 & pi0231;
assign w10010 = ~w9926 & ~pi0515;
assign w10011 = w9927 & pi0206;
assign w10012 = ~w9926 & ~pi0516;
assign w10013 = w9927 & pi0195;
assign w10014 = ~w9926 & ~pi0517;
assign w10015 = w9927 & pi0191;
assign w10016 = ~w9914 & ~pi0519;
assign w10017 = ~w9914 & ~pi0520;
assign w10018 = w9915 & pi0951;
assign w10019 = ~w9914 & ~pi0521;
assign w10020 = w9915 & pi0916;
assign w10021 = ~w9914 & ~pi0522;
assign w10022 = w9915 & pi0870;
assign w10023 = ~w9914 & ~pi0523;
assign w10024 = w9915 & pi0818;
assign w10025 = ~w9914 & ~pi0524;
assign w10026 = w9915 & pi0481;
assign w10027 = ~w9914 & ~pi0525;
assign w10028 = w9915 & pi0231;
assign w10029 = ~w9914 & ~pi0526;
assign w10030 = w9915 & pi0211;
assign w10031 = ~w9914 & ~pi0527;
assign w10032 = w9915 & pi0206;
assign w10033 = ~w9914 & ~pi0528;
assign w10034 = w9915 & pi0191;
assign w10035 = ~w9908 & ~pi0530;
assign w10036 = ~w9908 & ~pi0531;
assign w10037 = w9909 & pi0950;
assign w10038 = ~w9908 & ~pi0532;
assign w10039 = w9909 & pi0915;
assign w10040 = ~w9908 & ~pi0533;
assign w10041 = w9909 & pi0882;
assign w10042 = ~w9908 & ~pi0534;
assign w10043 = w9909 & pi0866;
assign w10044 = ~w9908 & ~pi0535;
assign w10045 = w9909 & pi0479;
assign w10046 = ~w9908 & ~pi0536;
assign w10047 = w9909 & pi0334;
assign w10048 = ~w9908 & ~pi0537;
assign w10049 = w9909 & pi0235;
assign w10050 = ~w9908 & ~pi0538;
assign w10051 = w9909 & pi0207;
assign w10052 = ~w9908 & ~pi0539;
assign w10053 = w9909 & pi0196;
assign w10054 = ~w9908 & ~pi0540;
assign w10055 = w9909 & pi0192;
assign w10056 = ~w9906 & ~pi0542;
assign w10057 = ~w9948 & ~pi0543;
assign w10058 = ~w9948 & ~pi0544;
assign w10059 = w9948 & w3363;
assign w10060 = w10059 & pi0915;
assign w10061 = ~w9948 & ~pi0545;
assign w10062 = w10059 & pi0882;
assign w10063 = ~w9948 & ~pi0546;
assign w10064 = w10059 & pi0866;
assign w10065 = ~w9948 & ~pi0547;
assign w10066 = w10059 & pi0819;
assign w10067 = ~w9948 & ~pi0548;
assign w10068 = w10059 & pi0479;
assign w10069 = ~w9948 & ~pi0549;
assign w10070 = w10059 & pi0334;
assign w10071 = ~w9948 & ~pi0550;
assign w10072 = w10059 & pi0235;
assign w10073 = ~w9948 & ~pi0551;
assign w10074 = w10059 & pi0212;
assign w10075 = ~w9948 & ~pi0552;
assign w10076 = w10059 & pi0207;
assign w10077 = ~w9948 & ~pi0553;
assign w10078 = w10059 & pi0950;
assign w10079 = ~w9948 & ~pi0554;
assign w10080 = w10059 & pi0196;
assign w10081 = ~w9948 & ~pi0555;
assign w10082 = w10059 & pi0192;
assign w10083 = ~w9752 & ~pi0557;
assign w10084 = ~w9752 & ~pi0558;
assign w10085 = ~w9942 & ~pi0559;
assign w10086 = ~w9942 & ~pi0560;
assign w10087 = ~w9942 & ~pi0561;
assign w10088 = ~w9908 & ~pi0562;
assign w10089 = ~w9942 & ~pi0563;
assign w10090 = ~w9768 & ~pi0564;
assign w10091 = ~w9768 & ~pi0565;
assign w10092 = ~w9768 & ~pi0566;
assign w10093 = ~w9908 & ~pi0567;
assign w10094 = ~w9908 & ~pi0568;
assign w10095 = ~w9768 & ~pi0569;
assign w10096 = ~w9768 & ~pi0570;
assign w10097 = ~w9768 & ~pi0571;
assign w10098 = ~w9768 & ~pi0572;
assign w10099 = ~w9768 & ~pi0573;
assign w10100 = ~w9768 & ~pi0574;
assign w10101 = ~w9768 & ~pi0575;
assign w10102 = ~w9768 & ~pi0576;
assign w10103 = ~w9768 & ~pi0577;
assign w10104 = ~w9795 & ~pi0578;
assign w10105 = ~w9795 & ~pi0579;
assign w10106 = ~w9795 & ~pi0580;
assign w10107 = ~w9795 & ~pi0581;
assign w10108 = ~w9795 & ~pi0582;
assign w10109 = ~w9795 & ~pi0583;
assign w10110 = ~w9795 & ~pi0584;
assign w10111 = ~w9768 & ~pi0585;
assign w10112 = ~w9795 & ~pi0586;
assign w10113 = ~w9795 & ~pi0587;
assign w10114 = ~w9795 & ~pi0588;
assign w10115 = ~w9795 & ~pi0589;
assign w10116 = ~w9795 & ~pi0590;
assign w10117 = ~w9795 & ~pi0591;
assign w10118 = ~w9795 & ~pi0592;
assign w10119 = ~w9752 & ~pi0593;
assign w10120 = ~w9752 & ~pi0594;
assign w10121 = ~w9752 & ~pi0595;
assign w10122 = ~w9752 & ~pi0596;
assign w10123 = ~w9752 & ~pi0597;
assign w10124 = ~w9752 & ~pi0598;
assign w10125 = ~w9752 & ~pi0599;
assign w10126 = ~w9752 & ~pi0600;
assign w10127 = ~pi0601 & pi1036;
assign w10128 = ~w9906 & ~pi0603;
assign w10129 = ~w9765 & ~pi0604;
assign w10130 = ~w9906 & ~pi0605;
assign w10131 = ~w9906 & ~pi0606;
assign w10132 = ~w9765 & ~pi0607;
assign w10133 = w9765 & w2398;
assign w10134 = w10133 & pi0947;
assign w10135 = ~w9765 & ~pi0608;
assign w10136 = w10133 & pi0923;
assign w10137 = ~w9765 & ~pi0609;
assign w10138 = w10133 & pi0877;
assign w10139 = ~w9765 & ~pi0610;
assign w10140 = w10133 & pi0871;
assign w10141 = ~w9765 & ~pi0611;
assign w10142 = w10133 & pi0814;
assign w10143 = ~w9765 & ~pi0612;
assign w10144 = w10133 & pi0480;
assign w10145 = ~w9765 & ~pi0613;
assign w10146 = w9906 & w3363;
assign w10147 = w10146 & pi0915;
assign w10148 = ~w9906 & ~pi0614;
assign w10149 = w10133 & pi0335;
assign w10150 = ~w9765 & ~pi0615;
assign w10151 = w10133 & pi0233;
assign w10152 = ~w9765 & ~pi0616;
assign w10153 = w10146 & pi0882;
assign w10154 = ~w9906 & ~pi0617;
assign w10155 = w10133 & pi0213;
assign w10156 = ~w9765 & ~pi0618;
assign w10157 = w10133 & pi0208;
assign w10158 = ~w9765 & ~pi0619;
assign w10159 = ~w9765 & ~pi0620;
assign w10160 = w10133 & pi0197;
assign w10161 = ~w9765 & ~pi0621;
assign w10162 = w10133 & pi0193;
assign w10163 = ~w9765 & ~pi0623;
assign w10164 = w10146 & pi0479;
assign w10165 = ~w9906 & ~pi0624;
assign w10166 = ~w9765 & ~pi0625;
assign w10167 = w10146 & pi0334;
assign w10168 = ~w9906 & ~pi0626;
assign w10169 = w10146 & pi0235;
assign w10170 = ~w9906 & ~pi0627;
assign w10171 = ~w9765 & ~pi0628;
assign w10172 = w10146 & pi0212;
assign w10173 = ~w9906 & ~pi0629;
assign w10174 = ~w9765 & ~pi0630;
assign w10175 = ~w9765 & ~pi0631;
assign w10176 = w10146 & pi0207;
assign w10177 = ~w9906 & ~pi0632;
assign w10178 = ~w9765 & ~pi0633;
assign w10179 = ~w9906 & ~pi0634;
assign w10180 = w2398 & pi0635;
assign w10181 = ~w2398 & ~pi0635;
assign w10182 = ~pi1834 & pi2020;
assign w10183 = ~w9906 & ~pi0637;
assign w10184 = ~w9765 & ~pi0638;
assign w10185 = ~w9908 & ~pi0639;
assign w10186 = ~w9906 & ~pi0641;
assign w10187 = ~w9960 & ~pi0642;
assign w10188 = ~w9914 & ~pi0643;
assign w10189 = w9914 & pi0643;
assign w10190 = pi1145 & pi0643;
assign w10191 = pi1145 & ~w10188;
assign w10192 = ~w9960 & ~pi0644;
assign w10193 = ~w9948 & ~pi0645;
assign w10194 = ~w9960 & ~pi0646;
assign w10195 = w9960 & w3383;
assign w10196 = w10195 & pi0333;
assign w10197 = ~w9960 & ~pi0647;
assign w10198 = ~w9948 & ~pi0648;
assign w10199 = ~w9960 & ~pi0649;
assign w10200 = ~w9960 & ~pi0650;
assign w10201 = ~w9948 & ~pi0651;
assign w10202 = ~w9948 & ~pi0652;
assign w10203 = ~w9948 & ~pi0653;
assign w10204 = ~w9948 & ~pi0654;
assign w10205 = ~w9908 & ~pi0655;
assign w10206 = w10146 & pi0866;
assign w10207 = ~w9906 & ~pi0656;
assign w10208 = ~pi1834 & ~pi0635;
assign w10209 = ~w9926 & ~pi0658;
assign w10210 = ~w9908 & ~pi0659;
assign w10211 = ~w9908 & ~pi0660;
assign w10212 = ~w9914 & ~pi0661;
assign w10213 = ~w9914 & ~pi0662;
assign w10214 = ~w9914 & ~pi0663;
assign w10215 = ~w9926 & ~pi0664;
assign w10216 = ~w9926 & ~pi0665;
assign w10217 = ~w9948 & ~pi0666;
assign w10218 = ~w9942 & ~pi0667;
assign w10219 = ~w9942 & ~pi0668;
assign w10220 = ~w9942 & ~pi0669;
assign w10221 = ~w9942 & ~pi0670;
assign w10222 = ~w9942 & ~pi0671;
assign w10223 = ~w9942 & ~pi0672;
assign w10224 = ~w9942 & ~pi0673;
assign w10225 = ~w9942 & ~pi0674;
assign w10226 = ~w9934 & ~pi0675;
assign w10227 = ~w9934 & ~pi0676;
assign w10228 = ~w9934 & ~pi0677;
assign w10229 = ~w9934 & ~pi0678;
assign w10230 = ~w9934 & ~pi0679;
assign w10231 = ~w9934 & ~pi0680;
assign w10232 = ~w9934 & ~pi0681;
assign w10233 = ~w9934 & ~pi0682;
assign w10234 = ~w9934 & ~pi0683;
assign w10235 = ~w9934 & ~pi0684;
assign w10236 = ~w9934 & ~pi0685;
assign w10237 = ~w9934 & ~pi0686;
assign w10238 = ~w9934 & ~pi0687;
assign w10239 = ~w9934 & ~pi0688;
assign w10240 = ~w9934 & ~pi0689;
assign w10241 = ~w9926 & ~pi0690;
assign w10242 = ~w9926 & ~pi0691;
assign w10243 = ~w9926 & ~pi0692;
assign w10244 = ~w9926 & ~pi0693;
assign w10245 = ~w9926 & ~pi0694;
assign w10246 = ~w9926 & ~pi0695;
assign w10247 = ~w9926 & ~pi0696;
assign w10248 = ~w9926 & ~pi0697;
assign w10249 = ~w9942 & ~pi0698;
assign w10250 = ~w9926 & ~pi0699;
assign w10251 = ~w9942 & ~pi0700;
assign w10252 = ~w9926 & ~pi0701;
assign w10253 = ~w9926 & ~pi0702;
assign w10254 = ~w9926 & ~pi0703;
assign w10255 = ~w9926 & ~pi0704;
assign w10256 = ~w9914 & ~pi0705;
assign w10257 = ~w9914 & ~pi0706;
assign w10258 = ~w9914 & ~pi0707;
assign w10259 = ~w9914 & ~pi0708;
assign w10260 = ~w9914 & ~pi0709;
assign w10261 = ~w9914 & ~pi0710;
assign w10262 = ~w9926 & ~pi0711;
assign w10263 = ~w9914 & ~pi0712;
assign w10264 = ~w9914 & ~pi0713;
assign w10265 = ~w9942 & ~pi0714;
assign w10266 = ~w9914 & ~pi0715;
assign w10267 = ~w9914 & ~pi0716;
assign w10268 = ~w9914 & ~pi0717;
assign w10269 = ~w9914 & ~pi0718;
assign w10270 = ~w9914 & ~pi0719;
assign w10271 = ~w9942 & ~pi0720;
assign w10272 = ~w9914 & ~pi0721;
assign w10273 = ~w9914 & ~pi0722;
assign w10274 = ~w9908 & ~pi0723;
assign w10275 = ~w9908 & ~pi0724;
assign w10276 = ~w9908 & ~pi0725;
assign w10277 = ~w9908 & ~pi0726;
assign w10278 = ~w9908 & ~pi0727;
assign w10279 = ~w9908 & ~pi0728;
assign w10280 = ~w9908 & ~pi0729;
assign w10281 = ~w9908 & ~pi0730;
assign w10282 = ~w9908 & ~pi0731;
assign w10283 = ~w9908 & ~pi0732;
assign w10284 = ~w9908 & ~pi0733;
assign w10285 = ~w9948 & ~pi0734;
assign w10286 = ~w9948 & ~pi0735;
assign w10287 = ~w9948 & ~pi0736;
assign w10288 = ~w9948 & ~pi0737;
assign w10289 = ~w9948 & ~pi0738;
assign w10290 = ~w9934 & ~pi0739;
assign w10291 = ~w9948 & ~pi0740;
assign w10292 = ~w9948 & ~pi0741;
assign w10293 = ~w9948 & ~pi0742;
assign w10294 = ~w9948 & ~pi0743;
assign w10295 = ~w9942 & ~pi0744;
assign w10296 = ~w9948 & ~pi0745;
assign w10297 = ~w9914 & pi1145;
assign w10298 = ~w9934 & ~pi0747;
assign w10299 = ~w9934 & ~pi0748;
assign w10300 = ~w9942 & ~pi0749;
assign w10301 = w10146 & pi0819;
assign w10302 = ~w9906 & ~pi0750;
assign w10303 = ~w9906 & ~pi0752;
assign w10304 = ~w9906 & ~pi0753;
assign w10305 = ~w9960 & ~pi0754;
assign w10306 = ~w9960 & ~pi0755;
assign w10307 = ~w9960 & ~pi0756;
assign w10308 = ~w9960 & ~pi0757;
assign w10309 = ~w9960 & ~pi0758;
assign w10310 = ~w9960 & ~pi0759;
assign w10311 = ~w9960 & ~pi0760;
assign w10312 = ~w9960 & ~pi0761;
assign w10313 = w10195 & pi0951;
assign w10314 = ~w9960 & ~pi0762;
assign w10315 = w10195 & pi0916;
assign w10316 = ~w9960 & ~pi0763;
assign w10317 = w10195 & pi0883;
assign w10318 = ~w9960 & ~pi0764;
assign w10319 = w10195 & pi0870;
assign w10320 = ~w9960 & ~pi0765;
assign w10321 = w10195 & pi0818;
assign w10322 = ~w9960 & ~pi0766;
assign w10323 = w10195 & pi0481;
assign w10324 = ~w9960 & ~pi0767;
assign w10325 = w10195 & pi0231;
assign w10326 = ~w9960 & ~pi0768;
assign w10327 = w10195 & pi0211;
assign w10328 = ~w9960 & ~pi0769;
assign w10329 = w10195 & pi0206;
assign w10330 = ~w9960 & ~pi0770;
assign w10331 = w10195 & pi0195;
assign w10332 = ~w9960 & ~pi0771;
assign w10333 = w10195 & pi0191;
assign w10334 = ~w9960 & ~pi0773;
assign w10335 = ~w9960 & ~pi0774;
assign w10336 = ~w9960 & ~pi0775;
assign w10337 = ~w9960 & ~pi0776;
assign w10338 = ~w9960 & ~pi0777;
assign w10339 = ~w9906 & ~pi0778;
assign w10340 = ~w9906 & ~pi0779;
assign w10341 = ~w9906 & ~pi0780;
assign w10342 = ~w9906 & ~pi0781;
assign w10343 = ~w9906 & ~pi0782;
assign w10344 = ~w9906 & ~pi0783;
assign w10345 = w10146 & pi0192;
assign w10346 = ~w9906 & ~pi0784;
assign w10347 = ~w9906 & ~pi0785;
assign w10348 = w10146 & pi0196;
assign w10349 = ~w9906 & ~pi0786;
assign w10350 = ~w9906 & ~pi0787;
assign w10351 = ~w9906 & ~pi0788;
assign w10352 = ~w9906 & ~pi0789;
assign w10353 = w3363 & pi0790;
assign w10354 = ~w3363 & ~pi0790;
assign w10355 = ~w9926 & ~pi0805;
assign w10356 = ~pi1076 & ~pi1903;
assign w10357 = ~pi1077 & ~pi1908;
assign w10358 = ~pi1876 & pi2055;
assign w10359 = ~pi0809 & ~pi0810;
assign w10360 = w10146 & pi0950;
assign w10361 = ~pi1876 & ~pi0790;
assign w10362 = w3383 & pi0821;
assign w10363 = ~w3383 & ~pi0821;
assign w10364 = ~pi0843 & pi1145;
assign w10365 = pi1881 & ~pi0821;
assign w10366 = pi1881 & pi2033;
assign w10367 = ~w4887 & pi1878;
assign w10368 = pi0893 & pi0897;
assign w10369 = ~pi0896 & ~pi0892;
assign w10370 = pi0896 & pi0892;
assign w10371 = ~pi0893 & ~pi0897;
assign w10372 = ~pi2239 & pi1198;
assign w10373 = ~w4917 & pi0810;
assign w10374 = w4917 & pi2026;
assign w10375 = pi2239 & pi1153;
assign w10376 = pi2240 & pi2146;
assign w10377 = ~pi2239 & pi1172;
assign w10378 = ~pi2240 & pi1844;
assign w10379 = w4917 & pi2130;
assign w10380 = ~w4922 & ~w4940;
assign w10381 = pi0932 & ~pi0924;
assign w10382 = w4887 & pi0932;
assign w10383 = ~pi0933 & ~pi0926;
assign w10384 = pi0933 & pi0926;
assign w10385 = pi1878 & pi0926;
assign w10386 = pi1878 & ~w10383;
assign w10387 = ~pi0930 & pi1169;
assign w10388 = ~pi0943 & ~pi0931;
assign w10389 = pi0943 & pi0931;
assign w10390 = w4887 & ~w5085;
assign w10391 = ~pi0933 & pi1878;
assign w10392 = ~pi0940 & ~pi0934;
assign w10393 = pi0940 & pi0934;
assign w10394 = ~pi0941 & ~pi0935;
assign w10395 = pi0941 & pi0935;
assign w10396 = ~pi0930 & ~pi0936;
assign w10397 = pi0930 & pi0936;
assign w10398 = ~pi0944 & ~pi0937;
assign w10399 = pi0944 & pi0937;
assign w10400 = ~pi0941 & pi1164;
assign w10401 = ~pi0943 & pi1176;
assign w10402 = ~pi0942 & ~pi0945;
assign w10403 = pi0942 & pi0945;
assign w10404 = ~pi1938 & pi0952;
assign w10405 = pi1938 & pi2174;
assign w10406 = ~pi1938 & pi0953;
assign w10407 = pi1938 & pi2197;
assign w10408 = ~pi1938 & pi0954;
assign w10409 = pi1938 & pi2196;
assign w10410 = ~pi1938 & pi0955;
assign w10411 = pi1938 & pi2179;
assign w10412 = ~pi1938 & pi0956;
assign w10413 = pi1938 & pi2176;
assign w10414 = ~pi1938 & pi0957;
assign w10415 = pi1938 & pi2169;
assign w10416 = ~pi1938 & pi0958;
assign w10417 = pi1938 & pi2173;
assign w10418 = ~pi1938 & pi0959;
assign w10419 = pi1938 & pi2167;
assign w10420 = ~pi1938 & pi0960;
assign w10421 = pi1938 & pi2166;
assign w10422 = ~pi1938 & pi0961;
assign w10423 = pi1938 & pi2192;
assign w10424 = pi0930 & pi0962;
assign w10425 = ~pi0930 & pi2174;
assign w10426 = pi0930 & pi0963;
assign w10427 = ~pi0930 & pi2197;
assign w10428 = pi0930 & pi0964;
assign w10429 = ~pi0930 & pi2196;
assign w10430 = pi0930 & pi0965;
assign w10431 = ~pi0930 & pi2179;
assign w10432 = pi0930 & pi0966;
assign w10433 = ~pi0930 & pi2176;
assign w10434 = pi0930 & pi0967;
assign w10435 = ~pi0930 & pi2169;
assign w10436 = pi0930 & pi0968;
assign w10437 = ~pi0930 & pi2173;
assign w10438 = pi0930 & pi0969;
assign w10439 = ~pi0930 & pi2167;
assign w10440 = pi0930 & pi0970;
assign w10441 = ~pi0930 & pi2166;
assign w10442 = pi0930 & pi0971;
assign w10443 = ~pi0930 & pi2192;
assign w10444 = pi0943 & pi0972;
assign w10445 = ~pi0943 & pi2174;
assign w10446 = pi0943 & pi0973;
assign w10447 = ~pi0943 & pi2197;
assign w10448 = pi0943 & pi0974;
assign w10449 = ~pi0943 & pi2196;
assign w10450 = pi0943 & pi0975;
assign w10451 = ~pi0943 & pi2179;
assign w10452 = pi0943 & pi0976;
assign w10453 = ~pi0943 & pi2176;
assign w10454 = pi0943 & pi0977;
assign w10455 = ~pi0943 & pi2169;
assign w10456 = pi0943 & pi0978;
assign w10457 = ~pi0943 & pi2173;
assign w10458 = pi0943 & pi0979;
assign w10459 = ~pi0943 & pi2167;
assign w10460 = pi0943 & pi0980;
assign w10461 = ~pi0943 & pi2166;
assign w10462 = pi0943 & pi0981;
assign w10463 = ~pi0943 & pi2192;
assign w10464 = ~pi1940 & pi0982;
assign w10465 = pi1940 & pi2174;
assign w10466 = ~pi1940 & pi0983;
assign w10467 = pi1940 & pi2197;
assign w10468 = ~pi1940 & pi0984;
assign w10469 = pi1940 & pi2196;
assign w10470 = ~pi1940 & pi0985;
assign w10471 = pi1940 & pi2179;
assign w10472 = ~pi1940 & pi0986;
assign w10473 = pi1940 & pi2176;
assign w10474 = ~pi1940 & pi0987;
assign w10475 = pi1940 & pi2169;
assign w10476 = ~pi1940 & pi0988;
assign w10477 = pi1940 & pi2173;
assign w10478 = ~pi1940 & pi0989;
assign w10479 = pi1940 & pi2167;
assign w10480 = ~pi1940 & pi0990;
assign w10481 = pi1940 & pi2166;
assign w10482 = ~pi1940 & pi0991;
assign w10483 = pi1940 & pi2192;
assign w10484 = pi0941 & pi0992;
assign w10485 = ~pi0941 & pi2172;
assign w10486 = pi0941 & pi0993;
assign w10487 = ~pi0941 & pi2168;
assign w10488 = pi0941 & pi0994;
assign w10489 = ~pi0941 & pi2178;
assign w10490 = ~pi1941 & pi0995;
assign w10491 = pi1941 & pi2186;
assign w10492 = ~pi1941 & pi0996;
assign w10493 = pi1941 & pi2172;
assign w10494 = ~pi1941 & pi0997;
assign w10495 = pi1941 & pi2168;
assign w10496 = ~pi1941 & pi0998;
assign w10497 = pi1941 & pi2193;
assign w10498 = pi0941 & pi0999;
assign w10499 = ~pi0941 & pi2198;
assign w10500 = pi0941 & pi1000;
assign w10501 = ~pi0941 & pi2187;
assign w10502 = ~pi1941 & pi1001;
assign w10503 = pi1941 & pi2170;
assign w10504 = ~pi1941 & pi1002;
assign w10505 = pi1941 & pi2182;
assign w10506 = ~pi1941 & pi1003;
assign w10507 = pi1941 & pi2175;
assign w10508 = ~pi1941 & pi1004;
assign w10509 = pi1941 & pi2177;
assign w10510 = pi0941 & pi1005;
assign w10511 = ~pi0941 & pi2181;
assign w10512 = ~pi1941 & pi1006;
assign w10513 = pi1941 & pi2167;
assign w10514 = ~pi1941 & pi1007;
assign w10515 = pi1941 & pi2188;
assign w10516 = pi0941 & pi1008;
assign w10517 = ~pi0941 & pi2191;
assign w10518 = pi0941 & pi1009;
assign w10519 = ~pi0941 & pi2175;
assign w10520 = pi0941 & pi1010;
assign w10521 = ~pi0941 & pi2184;
assign w10522 = pi0941 & pi1011;
assign w10523 = ~pi0941 & pi2188;
assign w10524 = pi2240 & ~pi1989;
assign w10525 = pi0941 & pi1013;
assign w10526 = ~pi0941 & pi2193;
assign w10527 = pi0940 & pi1941;
assign w10528 = ~pi1940 & pi1015;
assign w10529 = pi1940 & pi2185;
assign w10530 = pi0942 & pi1938;
assign w10531 = pi0930 & pi1019;
assign w10532 = ~pi0930 & pi2170;
assign w10533 = ~pi2239 & ~pi1989;
assign w10534 = pi0930 & pi1021;
assign w10535 = pi0930 & pi1022;
assign w10536 = ~pi0930 & pi2178;
assign w10537 = pi0930 & pi1023;
assign w10538 = pi0930 & pi1024;
assign w10539 = ~pi0930 & pi2172;
assign w10540 = pi0941 & pi1025;
assign w10541 = ~pi0941 & pi2176;
assign w10542 = ~pi0942 & pi1027;
assign w10543 = pi0942 & pi2192;
assign w10544 = ~pi0942 & pi1028;
assign w10545 = pi0942 & pi2188;
assign w10546 = ~pi0942 & pi1029;
assign w10547 = pi0942 & pi2177;
assign w10548 = ~pi1941 & pi1030;
assign w10549 = pi1941 & pi2178;
assign w10550 = pi0941 & pi1031;
assign w10551 = ~pi0941 & pi2196;
assign w10552 = ~pi0942 & pi1032;
assign w10553 = pi0942 & pi2171;
assign w10554 = ~pi0942 & pi1033;
assign w10555 = pi0942 & pi2181;
assign w10556 = pi0940 & pi1034;
assign w10557 = ~pi0940 & pi2184;
assign w10558 = pi2239 & ~pi1989;
assign w10559 = pi0941 & pi1038;
assign w10560 = ~pi0941 & pi2179;
assign w10561 = ~pi0942 & pi1040;
assign w10562 = pi0942 & pi2196;
assign w10563 = ~pi0942 & pi1041;
assign w10564 = pi0942 & pi2168;
assign w10565 = pi0941 & pi1043;
assign w10566 = ~pi1940 & pi1047;
assign w10567 = pi1940 & pi2177;
assign w10568 = ~pi0941 & pi1048;
assign w10569 = pi0941 & pi2191;
assign w10570 = pi0940 & pi1049;
assign w10571 = ~pi0940 & pi2187;
assign w10572 = pi0941 & pi1050;
assign w10573 = pi0940 & pi1051;
assign w10574 = ~pi0940 & pi2194;
assign w10575 = pi0942 & pi1053;
assign w10576 = ~pi0942 & pi2177;
assign w10577 = pi0942 & pi1054;
assign w10578 = ~pi0942 & pi2192;
assign w10579 = pi0942 & pi1055;
assign w10580 = ~pi0942 & pi2188;
assign w10581 = pi0942 & pi1056;
assign w10582 = ~pi0942 & pi2181;
assign w10583 = pi0940 & pi1057;
assign w10584 = ~pi0940 & pi2182;
assign w10585 = pi0941 & pi1058;
assign w10586 = ~pi0941 & pi2174;
assign w10587 = pi0940 & pi1059;
assign w10588 = ~pi0940 & pi2190;
assign w10589 = pi0942 & pi1060;
assign w10590 = ~pi0942 & pi2171;
assign w10591 = pi0942 & pi1061;
assign w10592 = ~pi0942 & pi2196;
assign w10593 = ~pi1940 & pi1062;
assign w10594 = pi1940 & pi2184;
assign w10595 = pi0944 & pi1063;
assign w10596 = ~pi0944 & pi2190;
assign w10597 = ~pi0941 & pi1064;
assign w10598 = pi0941 & pi2194;
assign w10599 = pi0942 & pi1065;
assign w10600 = ~pi0942 & pi2168;
assign w10601 = ~pi0944 & pi1066;
assign w10602 = pi0944 & pi2194;
assign w10603 = pi0940 & pi1067;
assign w10604 = ~pi0940 & pi2197;
assign w10605 = pi0940 & pi1068;
assign w10606 = ~pi0940 & pi2189;
assign w10607 = ~pi0941 & pi1069;
assign w10608 = pi0941 & pi2184;
assign w10609 = ~pi0941 & pi1070;
assign w10610 = pi0941 & pi2176;
assign w10611 = ~pi0941 & pi1071;
assign w10612 = pi0941 & pi2177;
assign w10613 = ~pi0941 & pi1072;
assign w10614 = pi0941 & pi2181;
assign w10615 = ~pi1940 & pi1073;
assign w10616 = pi1940 & pi2171;
assign w10617 = ~pi0941 & pi1074;
assign w10618 = pi0941 & pi2179;
assign w10619 = pi0943 & pi1081;
assign w10620 = ~pi0943 & pi2168;
assign w10621 = pi0940 & pi1082;
assign w10622 = ~pi0940 & pi2183;
assign w10623 = ~pi0944 & pi1083;
assign w10624 = pi0944 & pi2166;
assign w10625 = ~pi0941 & pi1084;
assign w10626 = pi0941 & pi2178;
assign w10627 = ~pi0941 & pi1085;
assign w10628 = pi0941 & pi2172;
assign w10629 = ~pi0941 & pi1086;
assign w10630 = pi0941 & pi2195;
assign w10631 = ~pi1940 & pi1087;
assign w10632 = pi1940 & pi2168;
assign w10633 = ~pi0944 & pi1088;
assign w10634 = pi0944 & pi2197;
assign w10635 = ~pi0944 & pi1089;
assign w10636 = pi0944 & pi2190;
assign w10637 = ~pi0944 & pi1090;
assign w10638 = pi0944 & pi2175;
assign w10639 = ~pi0941 & pi1091;
assign w10640 = pi0941 & pi2170;
assign w10641 = ~pi0941 & pi1092;
assign w10642 = ~pi0941 & pi1093;
assign w10643 = pi0941 & pi2189;
assign w10644 = ~pi0940 & pi1094;
assign w10645 = pi0940 & pi2195;
assign w10646 = ~pi0940 & pi1095;
assign w10647 = pi0940 & pi2184;
assign w10648 = ~pi0944 & pi1096;
assign w10649 = pi0944 & pi2187;
assign w10650 = ~pi0944 & pi1097;
assign w10651 = pi0944 & pi2189;
assign w10652 = ~pi0940 & pi1098;
assign w10653 = pi0940 & pi2194;
assign w10654 = ~pi0941 & pi1099;
assign w10655 = ~pi0940 & pi1100;
assign w10656 = pi0940 & pi2182;
assign w10657 = ~pi1940 & pi1101;
assign w10658 = pi1940 & pi2193;
assign w10659 = ~pi1940 & pi1102;
assign w10660 = pi1940 & pi2186;
assign w10661 = ~pi0940 & pi1103;
assign w10662 = pi0940 & pi2176;
assign w10663 = ~pi0940 & pi1104;
assign w10664 = pi0940 & pi2190;
assign w10665 = pi0944 & pi1940;
assign w10666 = ~pi0944 & pi1107;
assign w10667 = pi0944 & pi2183;
assign w10668 = ~pi0940 & pi1108;
assign w10669 = pi0940 & pi2189;
assign w10670 = pi0941 & pi1109;
assign w10671 = ~pi0941 & pi2194;
assign w10672 = ~pi0940 & pi1110;
assign w10673 = pi0940 & pi2178;
assign w10674 = ~pi0940 & pi1111;
assign w10675 = pi0940 & pi2183;
assign w10676 = pi0941 & pi1114;
assign w10677 = pi0943 & pi1117;
assign w10678 = ~pi0943 & pi2177;
assign w10679 = pi0943 & pi1118;
assign w10680 = ~pi0943 & pi2184;
assign w10681 = pi0943 & pi1122;
assign w10682 = ~pi0943 & pi2182;
assign w10683 = pi0944 & pi1123;
assign w10684 = ~pi0944 & pi2166;
assign w10685 = ~pi0943 & pi1124;
assign w10686 = pi0943 & pi2195;
assign w10687 = pi0944 & pi1127;
assign w10688 = ~pi0944 & pi2194;
assign w10689 = pi0944 & pi1135;
assign w10690 = ~pi0944 & pi2175;
assign w10691 = pi0943 & pi1136;
assign w10692 = ~pi0943 & pi2171;
assign w10693 = pi0941 & pi1225;
assign w10694 = ~pi0941 & pi2182;
assign w10695 = pi0941 & pi1227;
assign w10696 = ~pi0940 & pi1231;
assign w10697 = pi0940 & pi2186;
assign w10698 = pi0941 & pi1232;
assign w10699 = ~pi0941 & pi2177;
assign w10700 = ~pi0940 & pi1233;
assign w10701 = pi0940 & pi2172;
assign w10702 = pi0941 & pi1234;
assign w10703 = ~pi0941 & pi2173;
assign w10704 = ~pi0940 & pi1235;
assign w10705 = pi0940 & pi2168;
assign w10706 = ~pi0940 & pi1236;
assign w10707 = pi0940 & pi2174;
assign w10708 = pi0941 & pi1237;
assign w10709 = ~pi0941 & pi2167;
assign w10710 = ~pi0940 & pi1238;
assign w10711 = pi0940 & pi2197;
assign w10712 = ~pi0940 & pi1239;
assign w10713 = pi0940 & pi2196;
assign w10714 = ~pi0940 & pi1240;
assign w10715 = pi0940 & pi2193;
assign w10716 = pi0941 & pi1241;
assign w10717 = ~pi0940 & pi1242;
assign w10718 = pi0940 & pi2179;
assign w10719 = pi0941 & pi1243;
assign w10720 = ~pi0940 & pi1244;
assign w10721 = pi0940 & pi2198;
assign w10722 = pi0941 & pi1245;
assign w10723 = ~pi0941 & pi2166;
assign w10724 = ~pi0940 & pi1246;
assign w10725 = pi0940 & pi2185;
assign w10726 = ~pi0940 & pi1247;
assign w10727 = pi0940 & pi2187;
assign w10728 = pi0941 & pi1248;
assign w10729 = ~pi0941 & pi2195;
assign w10730 = ~pi0940 & pi1249;
assign w10731 = pi0940 & pi2171;
assign w10732 = ~pi0940 & pi1250;
assign w10733 = pi0940 & pi2169;
assign w10734 = pi0941 & pi1251;
assign w10735 = ~pi0941 & pi2192;
assign w10736 = ~pi0940 & pi1252;
assign w10737 = pi0940 & pi2170;
assign w10738 = ~pi0941 & pi1253;
assign w10739 = pi0941 & pi2186;
assign w10740 = ~pi0940 & pi1254;
assign w10741 = w4887 & pi1990;
assign w10742 = pi2003 & pi2001;
assign w10743 = ~pi1997 & ~pi1998;
assign w10744 = pi2000 & pi1999;
assign one = 1;
assign po0000 = pi1858;
assign po0001 = pi0898;
assign po0002 = pi1869;
assign po0003 = pi1867;
assign po0004 = pi1835;
assign po0005 = pi1866;
assign po0006 = pi1836;
assign po0007 = pi1864;
assign po0008 = pi1868;
assign po0009 = pi1863;
assign po0010 = pi1837;
assign po0011 = pi1862;
assign po0012 = pi1861;
assign po0013 = pi1860;
assign po0014 = pi1859;
assign po0015 = pi1865;
assign po0016 = pi1890;
assign po0017 = pi1893;
assign po0018 = pi1902;
assign po0019 = pi1892;
assign po0020 = pi1891;
assign po0021 = pi1889;
assign po0022 = pi1888;
assign po0023 = pi1887;
assign po0024 = pi1894;
assign po0025 = pi1900;
assign po0026 = pi1898;
assign po0027 = pi1897;
assign po0028 = pi1896;
assign po0029 = pi1899;
assign po0030 = pi1895;
assign po0031 = pi1882;
assign po0032 = pi1963;
assign po0033 = pi1945;
assign po0034 = pi2134;
assign po0035 = ~w0;
assign po0036 = pi0000;
assign po0037 = pi0924;
assign po0038 = pi0201;
assign po0039 = pi0198;
assign po0040 = pi0202;
assign po0041 = pi0199;
assign po0042 = pi0203;
assign po0043 = pi0204;
assign po0044 = pi0347;
assign po0045 = pi0348;
assign po0046 = pi0332;
assign po0047 = pi2204;
assign po0048 = w10;
assign po0049 = ~w13;
assign po0050 = ~w16;
assign po0051 = ~w19;
assign po0052 = w21;
assign po0053 = w22;
assign po0054 = ~w25;
assign po0055 = ~w28;
assign po0056 = ~w31;
assign po0057 = ~w34;
assign po0058 = w35;
assign po0059 = w36;
assign po0060 = w37;
assign po0061 = w38;
assign po0062 = w39;
assign po0063 = w40;
assign po0064 = ~w43;
assign po0065 = ~w46;
assign po0066 = ~w49;
assign po0067 = ~w52;
assign po0068 = ~w55;
assign po0069 = ~w58;
assign po0070 = ~w61;
assign po0071 = ~w64;
assign po0072 = w65;
assign po0073 = w66;
assign po0074 = w67;
assign po0075 = w68;
assign po0076 = w69;
assign po0077 = w70;
assign po0078 = w71;
assign po0079 = w72;
assign po0080 = w73;
assign po0081 = w74;
assign po0082 = w75;
assign po0083 = w76;
assign po0084 = ~w79;
assign po0085 = ~w82;
assign po0086 = ~w85;
assign po0087 = ~w88;
assign po0088 = ~w91;
assign po0089 = ~w94;
assign po0090 = ~w97;
assign po0091 = ~w100;
assign po0092 = ~w103;
assign po0093 = ~w106;
assign po0094 = ~w109;
assign po0095 = ~w112;
assign po0096 = ~w115;
assign po0097 = ~w118;
assign po0098 = ~w121;
assign po0099 = ~w124;
assign po0100 = w125;
assign po0101 = w126;
assign po0102 = w127;
assign po0103 = w128;
assign po0104 = ~w131;
assign po0105 = ~w134;
assign po0106 = ~w137;
assign po0107 = ~w140;
assign po0108 = ~w143;
assign po0109 = ~w146;
assign po0110 = ~w149;
assign po0111 = ~w152;
assign po0112 = ~w155;
assign po0113 = ~w158;
assign po0114 = ~w161;
assign po0115 = ~w164;
assign po0116 = ~w167;
assign po0117 = ~w170;
assign po0118 = ~w173;
assign po0119 = ~w176;
assign po0120 = ~w179;
assign po0121 = ~w182;
assign po0122 = ~w185;
assign po0123 = ~w188;
assign po0124 = ~w191;
assign po0125 = ~w194;
assign po0126 = ~w197;
assign po0127 = ~w200;
assign po0128 = ~w203;
assign po0129 = ~w206;
assign po0130 = ~w209;
assign po0131 = ~w212;
assign po0132 = ~w215;
assign po0133 = ~w218;
assign po0134 = ~w221;
assign po0135 = ~w224;
assign po0136 = ~w227;
assign po0137 = ~w230;
assign po0138 = ~w233;
assign po0139 = ~w236;
assign po0140 = ~w239;
assign po0141 = ~w242;
assign po0142 = ~w245;
assign po0143 = ~w248;
assign po0144 = w249;
assign po0145 = w250;
assign po0146 = w251;
assign po0147 = w252;
assign po0148 = w253;
assign po0149 = w254;
assign po0150 = w255;
assign po0151 = w256;
assign po0152 = w257;
assign po0153 = w258;
assign po0154 = w259;
assign po0155 = w260;
assign po0156 = w261;
assign po0157 = w262;
assign po0158 = w263;
assign po0159 = w264;
assign po0160 = w265;
assign po0161 = w266;
assign po0162 = w267;
assign po0163 = w268;
assign po0164 = ~w271;
assign po0165 = ~w274;
assign po0166 = ~w277;
assign po0167 = ~w280;
assign po0168 = ~w283;
assign po0169 = ~w286;
assign po0170 = ~w289;
assign po0171 = ~w292;
assign po0172 = ~w295;
assign po0173 = ~w298;
assign po0174 = ~w301;
assign po0175 = ~w304;
assign po0176 = ~w307;
assign po0177 = ~w310;
assign po0178 = ~w313;
assign po0179 = ~w316;
assign po0180 = ~w319;
assign po0181 = ~w322;
assign po0182 = ~w325;
assign po0183 = ~w328;
assign po0184 = ~w331;
assign po0185 = ~w334;
assign po0186 = ~w337;
assign po0187 = ~w340;
assign po0188 = ~w343;
assign po0189 = ~w346;
assign po0190 = ~w349;
assign po0191 = ~w352;
assign po0192 = ~w355;
assign po0193 = ~w358;
assign po0194 = ~w361;
assign po0195 = ~w364;
assign po0196 = ~w367;
assign po0197 = ~w370;
assign po0198 = ~w373;
assign po0199 = ~w376;
assign po0200 = ~w379;
assign po0201 = ~w382;
assign po0202 = ~w385;
assign po0203 = ~w388;
assign po0204 = ~w391;
assign po0205 = ~w394;
assign po0206 = ~w397;
assign po0207 = ~w400;
assign po0208 = ~w403;
assign po0209 = ~w406;
assign po0210 = ~w409;
assign po0211 = ~w412;
assign po0212 = ~w415;
assign po0213 = ~w418;
assign po0214 = ~w421;
assign po0215 = ~w424;
assign po0216 = ~w427;
assign po0217 = ~w430;
assign po0218 = ~w433;
assign po0219 = ~w436;
assign po0220 = ~w439;
assign po0221 = ~w442;
assign po0222 = ~w445;
assign po0223 = ~w448;
assign po0224 = ~w451;
assign po0225 = ~w454;
assign po0226 = ~w457;
assign po0227 = ~w460;
assign po0228 = ~w463;
assign po0229 = ~w466;
assign po0230 = ~w469;
assign po0231 = ~w472;
assign po0232 = ~w475;
assign po0233 = ~w478;
assign po0234 = ~w481;
assign po0235 = ~w484;
assign po0236 = ~w487;
assign po0237 = ~w490;
assign po0238 = ~w493;
assign po0239 = ~w496;
assign po0240 = ~w499;
assign po0241 = ~w502;
assign po0242 = ~w505;
assign po0243 = ~w508;
assign po0244 = ~w511;
assign po0245 = ~w514;
assign po0246 = pi2200;
assign po0247 = one;
assign po0248 = pi2199;
assign po0249 = w524;
assign po0250 = w534;
assign po0251 = ~w537;
assign po0252 = w547;
assign po0253 = w557;
assign po0254 = w567;
assign po0255 = w577;
assign po0256 = ~w580;
assign po0257 = ~w583;
assign po0258 = ~w586;
assign po0259 = ~w589;
assign po0260 = pi0228;
assign po0261 = ~w592;
assign po0262 = ~w595;
assign po0263 = ~w598;
assign po0264 = ~w601;
assign po0265 = w609;
assign po0266 = w620;
assign po0267 = w628;
assign po0268 = w636;
assign po0269 = w644;
assign po0270 = w652;
assign po0271 = w655;
assign po0272 = w658;
assign po0273 = w661;
assign po0274 = w664;
assign po0275 = w667;
assign po0276 = w670;
assign po0277 = w673;
assign po0278 = w676;
assign po0279 = pi0331;
assign po0280 = w687;
assign po0281 = w689;
assign po0282 = ~w692;
assign po0283 = ~w695;
assign po0284 = ~w698;
assign po0285 = ~w701;
assign po0286 = ~w704;
assign po0287 = w707;
assign po0288 = w710;
assign po0289 = w712;
assign po0290 = ~w717;
assign po0291 = ~w745;
assign po0292 = ~w763;
assign po0293 = ~w791;
assign po0294 = ~w809;
assign po0295 = ~w837;
assign po0296 = ~w855;
assign po0297 = ~w883;
assign po0298 = ~w901;
assign po0299 = w903;
assign po0300 = w905;
assign po0301 = w907;
assign po0302 = w909;
assign po0303 = ~w912;
assign po0304 = ~w915;
assign po0305 = ~w918;
assign po0306 = ~w921;
assign po0307 = ~w924;
assign po0308 = ~w927;
assign po0309 = ~w930;
assign po0310 = ~w933;
assign po0311 = ~w937;
assign po0312 = ~w941;
assign po0313 = w945;
assign po0314 = w949;
assign po0315 = ~w987;
assign po0316 = ~w1023;
assign po0317 = ~w1045;
assign po0318 = ~w1067;
assign po0319 = ~w1089;
assign po0320 = ~w1111;
assign po0321 = ~w1140;
assign po0322 = ~w1169;
assign po0323 = ~w1184;
assign po0324 = ~w1199;
assign po0325 = ~w1214;
assign po0326 = ~w1229;
assign po0327 = ~w1237;
assign po0328 = ~w1245;
assign po0329 = ~w1260;
assign po0330 = ~w1275;
assign po0331 = ~w1313;
assign po0332 = ~w1349;
assign po0333 = ~w1371;
assign po0334 = ~w1393;
assign po0335 = ~w1415;
assign po0336 = ~w1444;
assign po0337 = ~w1459;
assign po0338 = ~w1481;
assign po0339 = ~w1503;
assign po0340 = ~w1525;
assign po0341 = ~w1540;
assign po0342 = ~w1555;
assign po0343 = ~w1563;
assign po0344 = ~w1571;
assign po0345 = ~w1586;
assign po0346 = ~w1601;
assign po0347 = ~w1638;
assign po0348 = ~w1674;
assign po0349 = ~w1696;
assign po0350 = ~w1725;
assign po0351 = ~w1747;
assign po0352 = ~w1769;
assign po0353 = ~w1791;
assign po0354 = ~w1813;
assign po0355 = ~w1850;
assign po0356 = ~w1872;
assign po0357 = ~w1908;
assign po0358 = ~w1930;
assign po0359 = ~w1945;
assign po0360 = ~w1967;
assign po0361 = ~w1989;
assign po0362 = ~w2004;
assign po0363 = ~w2026;
assign po0364 = ~w2034;
assign po0365 = ~w2063;
assign po0366 = ~w2078;
assign po0367 = ~w2100;
assign po0368 = ~w2115;
assign po0369 = ~w2130;
assign po0370 = ~w2138;
assign po0371 = ~w2160;
assign po0372 = ~w2175;
assign po0373 = ~w2190;
assign po0374 = ~w2205;
assign po0375 = ~w2213;
assign po0376 = ~w2221;
assign po0377 = ~w2236;
assign po0378 = ~w2251;
assign po0379 = ~w2254;
assign po0380 = w2255;
assign po0381 = w2256;
assign po0382 = pi0456;
assign po0383 = w2266;
assign po0384 = ~w2269;
assign po0385 = ~w2272;
assign po0386 = ~w2275;
assign po0387 = ~w2278;
assign po0388 = ~w2306;
assign po0389 = ~w2332;
assign po0390 = ~w2350;
assign po0391 = ~w2368;
assign po0392 = w2369;
assign po0393 = w2370;
assign po0394 = w2371;
assign po0395 = w2372;
assign po0396 = ~w2397;
assign po0397 = w2406;
assign po0398 = w2416;
assign po0399 = w2426;
assign po0400 = ~w2429;
assign po0401 = ~w2432;
assign po0402 = ~w2435;
assign po0403 = ~w2438;
assign po0404 = ~w2440;
assign po0405 = ~w2444;
assign po0406 = ~w2452;
assign po0407 = ~w2458;
assign po0408 = ~w2462;
assign po0409 = ~w2465;
assign po0410 = ~w2468;
assign po0411 = ~w2471;
assign po0412 = ~w2474;
assign po0413 = ~w2477;
assign po0414 = ~w2480;
assign po0415 = ~w2483;
assign po0416 = ~w2486;
assign po0417 = ~w2489;
assign po0418 = ~w2492;
assign po0419 = ~w2495;
assign po0420 = ~w2498;
assign po0421 = ~w2501;
assign po0422 = ~w2505;
assign po0423 = ~w2508;
assign po0424 = ~w2511;
assign po0425 = ~w2514;
assign po0426 = ~w2517;
assign po0427 = ~w2520;
assign po0428 = ~w2523;
assign po0429 = ~w2526;
assign po0430 = ~w2529;
assign po0431 = ~w2532;
assign po0432 = ~w2535;
assign po0433 = ~w2538;
assign po0434 = ~w2541;
assign po0435 = ~w2544;
assign po0436 = ~w2547;
assign po0437 = ~w2550;
assign po0438 = ~w2553;
assign po0439 = ~w2556;
assign po0440 = ~w2559;
assign po0441 = ~w2562;
assign po0442 = ~w2565;
assign po0443 = ~w2568;
assign po0444 = ~w2571;
assign po0445 = ~w2574;
assign po0446 = ~w2577;
assign po0447 = ~w2580;
assign po0448 = ~w2583;
assign po0449 = ~w2586;
assign po0450 = ~w2595;
assign po0451 = ~w2603;
assign po0452 = ~w2611;
assign po0453 = ~w2619;
assign po0454 = ~w2627;
assign po0455 = ~w2635;
assign po0456 = ~w2638;
assign po0457 = ~w2646;
assign po0458 = ~w2649;
assign po0459 = ~w2652;
assign po0460 = ~w2660;
assign po0461 = ~w2668;
assign po0462 = w2671;
assign po0463 = w2674;
assign po0464 = ~w2710;
assign po0465 = ~w2746;
assign po0466 = ~w2775;
assign po0467 = ~w2797;
assign po0468 = ~w2812;
assign po0469 = ~w2834;
assign po0470 = ~w2856;
assign po0471 = ~w2871;
assign po0472 = ~w2900;
assign po0473 = ~w2915;
assign po0474 = ~w2930;
assign po0475 = ~w2938;
assign po0476 = ~w2946;
assign po0477 = ~w2961;
assign po0478 = ~w2976;
assign po0479 = ~w3013;
assign po0480 = ~w3049;
assign po0481 = ~w3071;
assign po0482 = ~w3093;
assign po0483 = ~w3122;
assign po0484 = ~w3144;
assign po0485 = ~w3166;
assign po0486 = ~w3195;
assign po0487 = ~w3210;
assign po0488 = ~w3225;
assign po0489 = ~w3233;
assign po0490 = ~w3248;
assign po0491 = ~w3263;
assign po0492 = ~w3271;
assign po0493 = ~w3279;
assign po0494 = ~w3287;
assign po0495 = ~w3290;
assign po0496 = ~w3293;
assign po0497 = ~w3301;
assign po0498 = ~w3309;
assign po0499 = ~w3312;
assign po0500 = ~w3316;
assign po0501 = ~w3318;
assign po0502 = ~w3320;
assign po0503 = ~w3322;
assign po0504 = ~w3324;
assign po0505 = ~w3332;
assign po0506 = ~w3347;
assign po0507 = pi0640;
assign po0508 = ~w3362;
assign po0509 = ~w3375;
assign po0510 = ~w3379;
assign po0511 = ~w3382;
assign po0512 = ~w3391;
assign po0513 = ~w3394;
assign po0514 = w3397;
assign po0515 = ~w3400;
assign po0516 = ~w3404;
assign po0517 = ~w3407;
assign po0518 = ~w3410;
assign po0519 = ~w3414;
assign po0520 = ~w3417;
assign po0521 = ~w3420;
assign po0522 = ~w3424;
assign po0523 = ~w3427;
assign po0524 = ~w3430;
assign po0525 = ~w3433;
assign po0526 = ~w3443;
assign po0527 = ~w3446;
assign po0528 = ~w3449;
assign po0529 = ~w3452;
assign po0530 = ~w3455;
assign po0531 = ~w3458;
assign po0532 = ~w3461;
assign po0533 = ~w3464;
assign po0534 = ~w3470;
assign po0535 = ~w3473;
assign po0536 = ~w3476;
assign po0537 = ~w3479;
assign po0538 = ~w3487;
assign po0539 = ~w3493;
assign po0540 = ~w3496;
assign po0541 = ~w3499;
assign po0542 = ~w3502;
assign po0543 = ~w3505;
assign po0544 = ~w3508;
assign po0545 = ~w3511;
assign po0546 = ~w3514;
assign po0547 = ~w3517;
assign po0548 = ~w3520;
assign po0549 = ~w3523;
assign po0550 = ~w3526;
assign po0551 = ~w3529;
assign po0552 = ~w3532;
assign po0553 = ~w3535;
assign po0554 = ~w3538;
assign po0555 = ~w3541;
assign po0556 = ~w3544;
assign po0557 = ~w3547;
assign po0558 = ~w3550;
assign po0559 = ~w3553;
assign po0560 = ~w3556;
assign po0561 = ~w3559;
assign po0562 = ~w3562;
assign po0563 = ~w3565;
assign po0564 = ~w3568;
assign po0565 = ~w3571;
assign po0566 = ~w3574;
assign po0567 = ~w3577;
assign po0568 = ~w3580;
assign po0569 = ~w3583;
assign po0570 = ~w3586;
assign po0571 = ~w3589;
assign po0572 = ~w3592;
assign po0573 = ~w3595;
assign po0574 = ~w3598;
assign po0575 = ~w3601;
assign po0576 = ~w3604;
assign po0577 = ~w3607;
assign po0578 = ~w3610;
assign po0579 = ~w3613;
assign po0580 = ~w3616;
assign po0581 = ~w3619;
assign po0582 = ~w3622;
assign po0583 = ~w3625;
assign po0584 = ~w3628;
assign po0585 = ~w3631;
assign po0586 = ~w3634;
assign po0587 = ~w3637;
assign po0588 = ~w3640;
assign po0589 = ~w3643;
assign po0590 = ~w3646;
assign po0591 = ~w3649;
assign po0592 = ~w3652;
assign po0593 = ~w3655;
assign po0594 = ~w3658;
assign po0595 = ~w3661;
assign po0596 = ~w3664;
assign po0597 = ~w3667;
assign po0598 = ~w3670;
assign po0599 = ~w3673;
assign po0600 = ~w3676;
assign po0601 = ~w3679;
assign po0602 = ~w3682;
assign po0603 = ~w3685;
assign po0604 = ~w3688;
assign po0605 = ~w3691;
assign po0606 = ~w3694;
assign po0607 = ~w3697;
assign po0608 = ~w3700;
assign po0609 = ~w3708;
assign po0610 = ~w3716;
assign po0611 = ~w3724;
assign po0612 = ~w3732;
assign po0613 = ~w3740;
assign po0614 = ~w3748;
assign po0615 = ~w3751;
assign po0616 = ~w3754;
assign po0617 = ~w3757;
assign po0618 = ~w3765;
assign po0619 = ~w3768;
assign po0620 = ~w3771;
assign po0621 = ~w3774;
assign po0622 = ~w3782;
assign po0623 = ~w3790;
assign po0624 = ~w3798;
assign po0625 = ~w3801;
assign po0626 = ~w3804;
assign po0627 = ~w3807;
assign po0628 = ~w3810;
assign po0629 = ~w3813;
assign po0630 = ~w3816;
assign po0631 = ~w3819;
assign po0632 = ~w3822;
assign po0633 = ~w3825;
assign po0634 = ~w3828;
assign po0635 = ~w3831;
assign po0636 = ~w3834;
assign po0637 = ~w3837;
assign po0638 = ~w3840;
assign po0639 = ~w3843;
assign po0640 = ~w3846;
assign po0641 = ~w3849;
assign po0642 = ~w3852;
assign po0643 = ~w3855;
assign po0644 = ~w3858;
assign po0645 = ~w3861;
assign po0646 = ~w3864;
assign po0647 = ~w3867;
assign po0648 = ~w3870;
assign po0649 = ~w3873;
assign po0650 = ~w3876;
assign po0651 = ~w3879;
assign po0652 = w3882;
assign po0653 = w3885;
assign po0654 = ~w3888;
assign po0655 = ~w3891;
assign po0656 = ~w3899;
assign po0657 = ~w3907;
assign po0658 = ~w3910;
assign po0659 = ~w3913;
assign po0660 = ~w3916;
assign po0661 = ~w3919;
assign po0662 = ~w3922;
assign po0663 = ~w3925;
assign po0664 = ~w3928;
assign po0665 = ~w3931;
assign po0666 = ~w3934;
assign po0667 = ~w3937;
assign po0668 = ~w3940;
assign po0669 = ~w3943;
assign po0670 = ~w3946;
assign po0671 = ~w3949;
assign po0672 = ~w3952;
assign po0673 = ~w3955;
assign po0674 = ~w3958;
assign po0675 = ~w3961;
assign po0676 = ~w3964;
assign po0677 = ~w3967;
assign po0678 = ~w3970;
assign po0679 = ~w3973;
assign po0680 = ~w3976;
assign po0681 = ~w3979;
assign po0682 = ~w3982;
assign po0683 = ~w3985;
assign po0684 = ~w3988;
assign po0685 = ~w3991;
assign po0686 = w3995;
assign po0687 = ~w3997;
assign po0688 = ~w4000;
assign po0689 = ~w4003;
assign po0690 = ~w4011;
assign po0691 = pi0840;
assign po0692 = ~w4019;
assign po0693 = ~w4028;
assign po0694 = w4031;
assign po0695 = ~w4039;
assign po0696 = ~w4047;
assign po0697 = ~w4055;
assign po0698 = ~w4058;
assign po0699 = ~w4061;
assign po0700 = ~w4069;
assign po0701 = ~w4077;
assign po0702 = ~w4080;
assign po0703 = ~w4088;
assign po0704 = ~w4091;
assign po0705 = ~w4099;
assign po0706 = ~w4102;
assign po0707 = ~w4105;
assign po0708 = ~w4109;
assign po0709 = ~w4117;
assign po0710 = ~w4120;
assign po0711 = ~w4123;
assign po0712 = ~w4126;
assign po0713 = ~w4134;
assign po0714 = ~w4142;
assign po0715 = ~w4150;
assign po0716 = ~w4153;
assign po0717 = ~w4156;
assign po0718 = ~w4159;
assign po0719 = ~w4162;
assign po0720 = ~w4165;
assign po0721 = ~w4168;
assign po0722 = ~w4176;
assign po0723 = ~w4179;
assign po0724 = ~w4187;
assign po0725 = ~w4190;
assign po0726 = ~w4198;
assign po0727 = ~w4206;
assign po0728 = ~w4209;
assign po0729 = ~w4212;
assign po0730 = ~w4220;
assign po0731 = ~w4228;
assign po0732 = ~w4231;
assign po0733 = ~w4234;
assign po0734 = ~w4237;
assign po0735 = ~w4245;
assign po0736 = ~w4248;
assign po0737 = ~w4251;
assign po0738 = ~w4259;
assign po0739 = ~w4267;
assign po0740 = ~w4270;
assign po0741 = ~w4273;
assign po0742 = ~w4276;
assign po0743 = ~w4284;
assign po0744 = ~w4287;
assign po0745 = ~w4290;
assign po0746 = ~w4293;
assign po0747 = ~w4296;
assign po0748 = ~w4299;
assign po0749 = ~w4302;
assign po0750 = ~w4305;
assign po0751 = ~w4313;
assign po0752 = ~w4316;
assign po0753 = ~w4319;
assign po0754 = ~w4322;
assign po0755 = ~w4325;
assign po0756 = ~w4328;
assign po0757 = ~w4331;
assign po0758 = ~w4334;
assign po0759 = ~w4337;
assign po0760 = ~w4340;
assign po0761 = ~w4343;
assign po0762 = ~w4346;
assign po0763 = ~w4349;
assign po0764 = ~w4352;
assign po0765 = ~w4360;
assign po0766 = ~w4363;
assign po0767 = ~w4366;
assign po0768 = ~w4369;
assign po0769 = ~w4372;
assign po0770 = ~w4375;
assign po0771 = ~w4378;
assign po0772 = ~w4386;
assign po0773 = ~w4389;
assign po0774 = ~w4392;
assign po0775 = ~w4395;
assign po0776 = ~w4398;
assign po0777 = ~w4401;
assign po0778 = ~w4404;
assign po0779 = ~w4407;
assign po0780 = ~w4410;
assign po0781 = ~w4413;
assign po0782 = ~w4416;
assign po0783 = ~w4419;
assign po0784 = ~w4422;
assign po0785 = ~w4425;
assign po0786 = ~w4428;
assign po0787 = ~w4431;
assign po0788 = ~w4434;
assign po0789 = ~w4437;
assign po0790 = ~w4440;
assign po0791 = ~w4443;
assign po0792 = ~w4446;
assign po0793 = ~w4449;
assign po0794 = ~w4452;
assign po0795 = ~w4455;
assign po0796 = ~w4458;
assign po0797 = w4461;
assign po0798 = ~w4464;
assign po0799 = ~w4467;
assign po0800 = ~w4470;
assign po0801 = ~w4473;
assign po0802 = ~w4476;
assign po0803 = ~w4479;
assign po0804 = ~w4482;
assign po0805 = ~w4485;
assign po0806 = ~w4488;
assign po0807 = ~w4491;
assign po0808 = ~w4494;
assign po0809 = ~w4497;
assign po0810 = ~w4500;
assign po0811 = ~w4503;
assign po0812 = ~w4506;
assign po0813 = ~w4509;
assign po0814 = ~w4512;
assign po0815 = ~w4515;
assign po0816 = ~w4518;
assign po0817 = ~w4521;
assign po0818 = ~w4524;
assign po0819 = ~w4527;
assign po0820 = ~w4530;
assign po0821 = ~w4533;
assign po0822 = ~w4536;
assign po0823 = ~w4539;
assign po0824 = ~w4542;
assign po0825 = ~w4545;
assign po0826 = ~w4548;
assign po0827 = ~w4551;
assign po0828 = ~w4554;
assign po0829 = ~w4557;
assign po0830 = ~w4560;
assign po0831 = ~w4563;
assign po0832 = ~w4566;
assign po0833 = ~w4569;
assign po0834 = ~w4572;
assign po0835 = ~w4575;
assign po0836 = ~w4578;
assign po0837 = ~w4581;
assign po0838 = ~w4584;
assign po0839 = ~w4587;
assign po0840 = ~w4590;
assign po0841 = w4594;
assign po0842 = ~w4597;
assign po0843 = ~w4600;
assign po0844 = ~w4603;
assign po0845 = ~w4606;
assign po0846 = ~w4609;
assign po0847 = ~w4612;
assign po0848 = ~w4615;
assign po0849 = ~w4618;
assign po0850 = ~w4621;
assign po0851 = ~w4624;
assign po0852 = ~w4627;
assign po0853 = ~w4630;
assign po0854 = ~w4633;
assign po0855 = ~w4636;
assign po0856 = ~w4639;
assign po0857 = ~w4641;
assign po0858 = ~w4643;
assign po0859 = ~w4645;
assign po0860 = ~w4649;
assign po0861 = w4651;
assign po0862 = ~w4654;
assign po0863 = ~w4657;
assign po0864 = ~w4661;
assign po0865 = ~w4664;
assign po0866 = w4666;
assign po0867 = ~w4669;
assign po0868 = ~w4672;
assign po0869 = ~w4675;
assign po0870 = ~w4678;
assign po0871 = ~w4681;
assign po0872 = w4685;
assign po0873 = ~w4688;
assign po0874 = ~w4691;
assign po0875 = ~w4694;
assign po0876 = ~w4697;
assign po0877 = ~w4700;
assign po0878 = ~w4703;
assign po0879 = ~w4706;
assign po0880 = ~w4709;
assign po0881 = ~w4712;
assign po0882 = ~w4715;
assign po0883 = ~w4718;
assign po0884 = ~w4721;
assign po0885 = ~w4724;
assign po0886 = ~w4727;
assign po0887 = w4729;
assign po0888 = ~w4733;
assign po0889 = w531;
assign po0890 = w521;
assign po0891 = pi0876;
assign po0892 = w4735;
assign po0893 = w4737;
assign po0894 = w4740;
assign po0895 = ~w4744;
assign po0896 = ~w4747;
assign po0897 = ~w4750;
assign po0898 = ~w4753;
assign po0899 = ~w4756;
assign po0900 = ~w4759;
assign po0901 = ~w4762;
assign po0902 = ~w4765;
assign po0903 = ~w4768;
assign po0904 = ~w4771;
assign po0905 = ~w4774;
assign po0906 = ~w4777;
assign po0907 = ~w4780;
assign po0908 = ~w4783;
assign po0909 = ~w4786;
assign po0910 = ~w4789;
assign po0911 = ~w4792;
assign po0912 = w564;
assign po0913 = w574;
assign po0914 = w544;
assign po0915 = w554;
assign po0916 = w4793;
assign po0917 = ~w4796;
assign po0918 = ~w4799;
assign po0919 = ~w4802;
assign po0920 = ~w4805;
assign po0921 = ~w4808;
assign po0922 = ~w4811;
assign po0923 = ~w4813;
assign po0924 = w4814;
assign po0925 = w4815;
assign po0926 = w4816;
assign po0927 = pi0891;
assign po0928 = ~w4819;
assign po0929 = ~w4822;
assign po0930 = ~w4829;
assign po0931 = w4835;
assign po0932 = ~w4838;
assign po0933 = ~w4841;
assign po0934 = ~w4844;
assign po0935 = ~w4851;
assign po0936 = ~w4858;
assign po0937 = ~w4865;
assign po0938 = ~w4872;
assign po0939 = ~w4879;
assign po0940 = w4883;
assign po0941 = ~w4886;
assign po0942 = pi0925;
assign po0943 = w4900;
assign po0944 = w4903;
assign po0945 = w4904;
assign po0946 = w4907;
assign po0947 = w4910;
assign po0948 = w4913;
assign po0949 = ~w4947;
assign po0950 = ~w4960;
assign po0951 = ~w4973;
assign po0952 = ~w4986;
assign po0953 = ~w4999;
assign po0954 = w5001;
assign po0955 = ~w5014;
assign po0956 = ~w5027;
assign po0957 = ~w5030;
assign po0958 = ~w5033;
assign po0959 = w2263;
assign po0960 = ~w5036;
assign po0961 = ~w5039;
assign po0962 = ~w5042;
assign po0963 = ~w5045;
assign po0964 = ~w5048;
assign po0965 = ~w5051;
assign po0966 = ~w5054;
assign po0967 = ~w5057;
assign po0968 = w5061;
assign po0969 = w5065;
assign po0970 = w5069;
assign po0971 = w5073;
assign po0972 = w5077;
assign po0973 = w5081;
assign po0974 = ~w5084;
assign po0975 = w5087;
assign po0976 = pi1768;
assign po0977 = w5091;
assign po0978 = w2413;
assign po0979 = w2423;
assign po0980 = ~w5098;
assign po0981 = w5103;
assign po0982 = w5109;
assign po0983 = w5113;
assign po0984 = w5116;
assign po0985 = w5121;
assign po0986 = w5127;
assign po0987 = w5131;
assign po0988 = w5136;
assign po0989 = ~w5143;
assign po0990 = ~w5150;
assign po0991 = w5154;
assign po0992 = w5157;
assign po0993 = w5161;
assign po0994 = w5164;
assign po0995 = w5168;
assign po0996 = w5173;
assign po0997 = pi1930;
assign po0998 = ~w5176;
assign po0999 = ~w5179;
assign po1000 = ~w5182;
assign po1001 = ~w5185;
assign po1002 = ~w5188;
assign po1003 = ~w5193;
assign po1004 = ~w5196;
assign po1005 = ~w5199;
assign po1006 = ~w5202;
assign po1007 = ~w5205;
assign po1008 = ~w5208;
assign po1009 = ~w5211;
assign po1010 = ~w5214;
assign po1011 = ~w5217;
assign po1012 = ~w5220;
assign po1013 = ~w5224;
assign po1014 = ~w5227;
assign po1015 = ~w5230;
assign po1016 = ~w5233;
assign po1017 = ~w5236;
assign po1018 = ~w5239;
assign po1019 = ~w5242;
assign po1020 = ~w5245;
assign po1021 = ~w5248;
assign po1022 = ~w5251;
assign po1023 = ~w5255;
assign po1024 = ~w5258;
assign po1025 = ~w5261;
assign po1026 = ~w5264;
assign po1027 = ~w5267;
assign po1028 = ~w5270;
assign po1029 = ~w5273;
assign po1030 = ~w5276;
assign po1031 = ~w5279;
assign po1032 = ~w5282;
assign po1033 = ~w5287;
assign po1034 = ~w5290;
assign po1035 = ~w5293;
assign po1036 = ~w5296;
assign po1037 = ~w5299;
assign po1038 = ~w5302;
assign po1039 = ~w5305;
assign po1040 = ~w5308;
assign po1041 = ~w5311;
assign po1042 = ~w5314;
assign po1043 = ~w5318;
assign po1044 = ~w5321;
assign po1045 = ~w5324;
assign po1046 = ~w5329;
assign po1047 = ~w5332;
assign po1048 = ~w5335;
assign po1049 = ~w5338;
assign po1050 = ~w5341;
assign po1051 = ~w5344;
assign po1052 = ~w5347;
assign po1053 = ~w5350;
assign po1054 = ~w5353;
assign po1055 = ~w5356;
assign po1056 = ~w5359;
assign po1057 = ~w5362;
assign po1058 = ~w5365;
assign po1059 = ~w5368;
assign po1060 = ~w5371;
assign po1061 = ~w5374;
assign po1062 = ~w5377;
assign po1063 = ~w5381;
assign po1064 = ~w5384;
assign po1065 = ~w5388;
assign po1066 = ~w5391;
assign po1067 = ~w5394;
assign po1068 = ~w5397;
assign po1069 = ~w5401;
assign po1070 = ~w5405;
assign po1071 = ~w5409;
assign po1072 = ~w5412;
assign po1073 = ~w5415;
assign po1074 = ~w5418;
assign po1075 = ~w5421;
assign po1076 = ~w5425;
assign po1077 = ~w5428;
assign po1078 = ~w5431;
assign po1079 = ~w5434;
assign po1080 = ~w5437;
assign po1081 = ~w5440;
assign po1082 = ~w5443;
assign po1083 = ~w5446;
assign po1084 = ~w5449;
assign po1085 = ~w5452;
assign po1086 = ~w5455;
assign po1087 = ~w5459;
assign po1088 = ~w5462;
assign po1089 = ~w5465;
assign po1090 = ~w5468;
assign po1091 = ~w5471;
assign po1092 = ~w5474;
assign po1093 = ~w5477;
assign po1094 = ~w5480;
assign po1095 = ~w5483;
assign po1096 = ~w5486;
assign po1097 = ~w5489;
assign po1098 = ~w5492;
assign po1099 = ~w5496;
assign po1100 = ~w5499;
assign po1101 = ~w5502;
assign po1102 = ~w5505;
assign po1103 = ~w5508;
assign po1104 = ~w5511;
assign po1105 = ~w5514;
assign po1106 = ~w5517;
assign po1107 = ~w5520;
assign po1108 = ~w5523;
assign po1109 = ~w5526;
assign po1110 = ~w5529;
assign po1111 = ~w5532;
assign po1112 = ~w5535;
assign po1113 = ~w5538;
assign po1114 = ~w5541;
assign po1115 = ~w5544;
assign po1116 = ~w5547;
assign po1117 = ~w5550;
assign po1118 = ~w5553;
assign po1119 = ~w5556;
assign po1120 = ~w5559;
assign po1121 = ~w5562;
assign po1122 = ~w5565;
assign po1123 = ~w5568;
assign po1124 = ~w5571;
assign po1125 = ~w5574;
assign po1126 = w629;
assign po1127 = w602;
assign po1128 = w613;
assign po1129 = w637;
assign po1130 = w645;
assign po1131 = w621;
assign po1132 = ~w5577;
assign po1133 = ~w5580;
assign po1134 = ~w5583;
assign po1135 = ~w5586;
assign po1136 = ~w5589;
assign po1137 = ~w5592;
assign po1138 = ~w5595;
assign po1139 = ~w5598;
assign po1140 = ~w5601;
assign po1141 = ~w5604;
assign po1142 = ~w5607;
assign po1143 = ~w5610;
assign po1144 = ~w5613;
assign po1145 = ~w5616;
assign po1146 = ~w5619;
assign po1147 = ~w5622;
assign po1148 = ~w5625;
assign po1149 = ~w5628;
assign po1150 = ~w5631;
assign po1151 = ~w5634;
assign po1152 = ~w5637;
assign po1153 = ~w5640;
assign po1154 = ~w5643;
assign po1155 = ~w5646;
assign po1156 = ~w5650;
assign po1157 = ~w5653;
assign po1158 = ~w5656;
assign po1159 = ~w5659;
assign po1160 = ~w5662;
assign po1161 = ~w5665;
assign po1162 = ~w5668;
assign po1163 = ~w5671;
assign po1164 = ~w5674;
assign po1165 = ~w5677;
assign po1166 = ~w5680;
assign po1167 = ~w5683;
assign po1168 = ~w5686;
assign po1169 = ~w5689;
assign po1170 = ~w5692;
assign po1171 = ~w5695;
assign po1172 = ~w5698;
assign po1173 = ~w5701;
assign po1174 = ~w5704;
assign po1175 = ~w5707;
assign po1176 = w5710;
assign po1177 = w5713;
assign po1178 = ~w5716;
assign po1179 = ~w5719;
assign po1180 = w5722;
assign po1181 = ~w5725;
assign po1182 = ~w5728;
assign po1183 = ~w5732;
assign po1184 = ~w5735;
assign po1185 = ~w5738;
assign po1186 = ~w5741;
assign po1187 = ~w5744;
assign po1188 = ~w5747;
assign po1189 = ~w5750;
assign po1190 = ~w5753;
assign po1191 = ~w5756;
assign po1192 = ~w5759;
assign po1193 = ~w5762;
assign po1194 = ~w5765;
assign po1195 = ~w5768;
assign po1196 = ~w5771;
assign po1197 = ~w5774;
assign po1198 = ~w5777;
assign po1199 = ~w5780;
assign po1200 = ~w5783;
assign po1201 = ~w5786;
assign po1202 = ~w5789;
assign po1203 = ~w5792;
assign po1204 = ~w5795;
assign po1205 = ~w5798;
assign po1206 = ~w5801;
assign po1207 = ~w5804;
assign po1208 = ~w5807;
assign po1209 = ~w5810;
assign po1210 = ~w5813;
assign po1211 = ~w5816;
assign po1212 = ~w5819;
assign po1213 = ~w5822;
assign po1214 = ~w5825;
assign po1215 = ~w5828;
assign po1216 = ~w5831;
assign po1217 = ~w5834;
assign po1218 = ~w5837;
assign po1219 = ~w5840;
assign po1220 = ~w5843;
assign po1221 = ~w5846;
assign po1222 = ~w5849;
assign po1223 = ~w5852;
assign po1224 = ~w5855;
assign po1225 = ~w5858;
assign po1226 = ~w5861;
assign po1227 = ~w5864;
assign po1228 = ~w5867;
assign po1229 = ~w5870;
assign po1230 = ~w5873;
assign po1231 = ~w5876;
assign po1232 = ~w5879;
assign po1233 = ~w5882;
assign po1234 = ~w5885;
assign po1235 = ~w5888;
assign po1236 = ~w5891;
assign po1237 = ~w5894;
assign po1238 = ~w5897;
assign po1239 = ~w5900;
assign po1240 = ~w5903;
assign po1241 = ~w5906;
assign po1242 = ~w5909;
assign po1243 = ~w5912;
assign po1244 = ~w5915;
assign po1245 = ~w5918;
assign po1246 = ~w5921;
assign po1247 = ~w5924;
assign po1248 = ~w5927;
assign po1249 = ~w5930;
assign po1250 = ~w5933;
assign po1251 = ~w5936;
assign po1252 = ~w5939;
assign po1253 = ~w5942;
assign po1254 = ~w5945;
assign po1255 = ~w5948;
assign po1256 = ~w5951;
assign po1257 = ~w5954;
assign po1258 = ~w5957;
assign po1259 = ~w5960;
assign po1260 = ~w5963;
assign po1261 = ~w5966;
assign po1262 = ~w5969;
assign po1263 = w5972;
assign po1264 = w5975;
assign po1265 = w5978;
assign po1266 = w5981;
assign po1267 = w5984;
assign po1268 = w5987;
assign po1269 = w5990;
assign po1270 = w5993;
assign po1271 = w5996;
assign po1272 = w5999;
assign po1273 = w6002;
assign po1274 = w6005;
assign po1275 = ~w6008;
assign po1276 = ~w6011;
assign po1277 = ~w6014;
assign po1278 = ~w6017;
assign po1279 = ~w6020;
assign po1280 = ~w6023;
assign po1281 = ~w6026;
assign po1282 = ~w6029;
assign po1283 = ~w6032;
assign po1284 = ~w6035;
assign po1285 = ~w6038;
assign po1286 = ~w6041;
assign po1287 = ~w6044;
assign po1288 = ~w6047;
assign po1289 = ~w6050;
assign po1290 = ~w6053;
assign po1291 = ~w6056;
assign po1292 = ~w6059;
assign po1293 = ~w6062;
assign po1294 = ~w6065;
assign po1295 = ~w6068;
assign po1296 = ~w6071;
assign po1297 = ~w6074;
assign po1298 = ~w6077;
assign po1299 = ~w6080;
assign po1300 = ~w6083;
assign po1301 = ~w6086;
assign po1302 = ~w6089;
assign po1303 = ~w6092;
assign po1304 = ~w6095;
assign po1305 = ~w6098;
assign po1306 = ~w6101;
assign po1307 = ~w6104;
assign po1308 = ~w6107;
assign po1309 = ~w6110;
assign po1310 = ~w6113;
assign po1311 = ~w6116;
assign po1312 = ~w6119;
assign po1313 = ~w6122;
assign po1314 = ~w6125;
assign po1315 = ~w6128;
assign po1316 = ~w6131;
assign po1317 = ~w6134;
assign po1318 = ~w6137;
assign po1319 = ~w6140;
assign po1320 = ~w6143;
assign po1321 = ~w6146;
assign po1322 = ~w6149;
assign po1323 = ~w6152;
assign po1324 = ~w6155;
assign po1325 = ~w6158;
assign po1326 = ~w6161;
assign po1327 = ~w6164;
assign po1328 = ~w6167;
assign po1329 = ~w6170;
assign po1330 = ~w6173;
assign po1331 = ~w6176;
assign po1332 = ~w6179;
assign po1333 = ~w6182;
assign po1334 = ~w6185;
assign po1335 = ~w6188;
assign po1336 = ~w6191;
assign po1337 = ~w6194;
assign po1338 = ~w6197;
assign po1339 = ~w6200;
assign po1340 = ~w6203;
assign po1341 = ~w6206;
assign po1342 = ~w6209;
assign po1343 = ~w6212;
assign po1344 = ~w6215;
assign po1345 = ~w6218;
assign po1346 = ~w6221;
assign po1347 = ~w6224;
assign po1348 = ~w6227;
assign po1349 = ~w6230;
assign po1350 = ~w6233;
assign po1351 = ~w6236;
assign po1352 = ~w6239;
assign po1353 = ~w6242;
assign po1354 = ~w6245;
assign po1355 = ~w6248;
assign po1356 = ~w6251;
assign po1357 = ~w6254;
assign po1358 = ~w6257;
assign po1359 = ~w6260;
assign po1360 = ~w6263;
assign po1361 = ~w6266;
assign po1362 = ~w6269;
assign po1363 = ~w6272;
assign po1364 = ~w6275;
assign po1365 = ~w6278;
assign po1366 = ~w6281;
assign po1367 = ~w6284;
assign po1368 = ~w6287;
assign po1369 = ~w6290;
assign po1370 = ~w6293;
assign po1371 = ~w6296;
assign po1372 = ~w6299;
assign po1373 = ~w6302;
assign po1374 = ~w6305;
assign po1375 = ~w6308;
assign po1376 = ~w6311;
assign po1377 = ~w6314;
assign po1378 = ~w6317;
assign po1379 = ~w6320;
assign po1380 = ~w6323;
assign po1381 = ~w6326;
assign po1382 = ~w6329;
assign po1383 = ~w6332;
assign po1384 = ~w6335;
assign po1385 = ~w6338;
assign po1386 = ~w6341;
assign po1387 = ~w6344;
assign po1388 = ~w6347;
assign po1389 = ~w6350;
assign po1390 = ~w6353;
assign po1391 = ~w6356;
assign po1392 = ~w6359;
assign po1393 = ~w6362;
assign po1394 = ~w6365;
assign po1395 = ~w6368;
assign po1396 = ~w6371;
assign po1397 = ~w6374;
assign po1398 = ~w6377;
assign po1399 = ~w6380;
assign po1400 = ~w6383;
assign po1401 = ~w6386;
assign po1402 = ~w6389;
assign po1403 = ~w6392;
assign po1404 = ~w6395;
assign po1405 = ~w6398;
assign po1406 = ~w6401;
assign po1407 = ~w6404;
assign po1408 = ~w6407;
assign po1409 = ~w6410;
assign po1410 = ~w6413;
assign po1411 = ~w6416;
assign po1412 = ~w6419;
assign po1413 = ~w6422;
assign po1414 = ~w6425;
assign po1415 = ~w6428;
assign po1416 = ~w6431;
assign po1417 = ~w6434;
assign po1418 = ~w6437;
assign po1419 = ~w6440;
assign po1420 = ~w6443;
assign po1421 = ~w6446;
assign po1422 = ~w6449;
assign po1423 = ~w6452;
assign po1424 = ~w6455;
assign po1425 = ~w6458;
assign po1426 = ~w6461;
assign po1427 = ~w6464;
assign po1428 = ~w6467;
assign po1429 = ~w6470;
assign po1430 = ~w6473;
assign po1431 = ~w6476;
assign po1432 = ~w6479;
assign po1433 = ~w6482;
assign po1434 = ~w6485;
assign po1435 = ~w6488;
assign po1436 = ~w6491;
assign po1437 = ~w6494;
assign po1438 = ~w6497;
assign po1439 = ~w6500;
assign po1440 = ~w6503;
assign po1441 = ~w6506;
assign po1442 = ~w6509;
assign po1443 = ~w6512;
assign po1444 = ~w6515;
assign po1445 = ~w6518;
assign po1446 = ~w6521;
assign po1447 = ~w6524;
assign po1448 = ~w6527;
assign po1449 = ~w6530;
assign po1450 = ~w6533;
assign po1451 = ~w6536;
assign po1452 = ~w6539;
assign po1453 = ~w6542;
assign po1454 = ~w6545;
assign po1455 = ~w6548;
assign po1456 = ~w6551;
assign po1457 = ~w6554;
assign po1458 = ~w6557;
assign po1459 = ~w6560;
assign po1460 = ~w6563;
assign po1461 = ~w6566;
assign po1462 = ~w6570;
assign po1463 = ~w6573;
assign po1464 = ~w6576;
assign po1465 = ~w6579;
assign po1466 = ~w6582;
assign po1467 = ~w6585;
assign po1468 = ~w6588;
assign po1469 = ~w6591;
assign po1470 = ~w6594;
assign po1471 = ~w6597;
assign po1472 = ~w6600;
assign po1473 = ~w6603;
assign po1474 = ~w6606;
assign po1475 = ~w6609;
assign po1476 = ~w6612;
assign po1477 = ~w6615;
assign po1478 = ~w6618;
assign po1479 = ~w6621;
assign po1480 = ~w6624;
assign po1481 = ~w6627;
assign po1482 = ~w6630;
assign po1483 = ~w6633;
assign po1484 = ~w6636;
assign po1485 = ~w6639;
assign po1486 = ~w6642;
assign po1487 = ~w6645;
assign po1488 = ~w6648;
assign po1489 = ~w6651;
assign po1490 = ~w6654;
assign po1491 = ~w6657;
assign po1492 = ~w6660;
assign po1493 = ~w6663;
assign po1494 = ~w6666;
assign po1495 = ~w6669;
assign po1496 = ~w6672;
assign po1497 = ~w6675;
assign po1498 = ~w6678;
assign po1499 = ~w6681;
assign po1500 = ~w6684;
assign po1501 = ~w6687;
assign po1502 = ~w6690;
assign po1503 = ~w6693;
assign po1504 = ~w6696;
assign po1505 = ~w6699;
assign po1506 = ~w6702;
assign po1507 = ~w6705;
assign po1508 = ~w6708;
assign po1509 = ~w6711;
assign po1510 = ~w6714;
assign po1511 = ~w6717;
assign po1512 = ~w6721;
assign po1513 = ~w6724;
assign po1514 = ~w6727;
assign po1515 = ~w6730;
assign po1516 = ~w6733;
assign po1517 = ~w6736;
assign po1518 = ~w6739;
assign po1519 = ~w6742;
assign po1520 = ~w6745;
assign po1521 = ~w6748;
assign po1522 = ~w6751;
assign po1523 = ~w6754;
assign po1524 = ~w6757;
assign po1525 = ~w6760;
assign po1526 = ~w6763;
assign po1527 = ~w6766;
assign po1528 = ~w6769;
assign po1529 = ~w6772;
assign po1530 = ~w6775;
assign po1531 = ~w6778;
assign po1532 = ~w6781;
assign po1533 = ~w6784;
assign po1534 = ~w6787;
assign po1535 = ~w6790;
assign po1536 = ~w6793;
assign po1537 = ~w6797;
assign po1538 = ~w6800;
assign po1539 = ~w6803;
assign po1540 = ~w6806;
assign po1541 = ~w6809;
assign po1542 = ~w6812;
assign po1543 = ~w6815;
assign po1544 = ~w6818;
assign po1545 = ~w6821;
assign po1546 = ~w6824;
assign po1547 = ~w6827;
assign po1548 = ~w6830;
assign po1549 = ~w6833;
assign po1550 = ~w6836;
assign po1551 = ~w6839;
assign po1552 = ~w6842;
assign po1553 = ~w6845;
assign po1554 = ~w6848;
assign po1555 = ~w6851;
assign po1556 = ~w6854;
assign po1557 = ~w6857;
assign po1558 = ~w6860;
assign po1559 = ~w6863;
assign po1560 = ~w6866;
assign po1561 = ~w6869;
assign po1562 = ~w6872;
assign po1563 = ~w6875;
assign po1564 = ~w6878;
assign po1565 = ~w6881;
assign po1566 = ~w6884;
assign po1567 = ~w6887;
assign po1568 = ~w6890;
assign po1569 = ~w6893;
assign po1570 = ~w6896;
assign po1571 = ~w6899;
assign po1572 = ~w6902;
assign po1573 = ~w6905;
assign po1574 = ~w6908;
assign po1575 = ~w6911;
assign po1576 = ~w6914;
assign po1577 = ~w6917;
assign po1578 = ~w6920;
assign po1579 = ~w6923;
assign po1580 = ~w6926;
assign po1581 = ~w6929;
assign po1582 = ~w6932;
assign po1583 = ~w6935;
assign po1584 = ~w6938;
assign po1585 = ~w6941;
assign po1586 = ~w6944;
assign po1587 = ~w6947;
assign po1588 = ~w6950;
assign po1589 = ~w6953;
assign po1590 = ~w6956;
assign po1591 = ~w6959;
assign po1592 = ~w6962;
assign po1593 = ~w6965;
assign po1594 = ~w6968;
assign po1595 = ~w6971;
assign po1596 = ~w6974;
assign po1597 = ~w6977;
assign po1598 = ~w6980;
assign po1599 = ~w6983;
assign po1600 = ~w6986;
assign po1601 = ~w6989;
assign po1602 = ~w6992;
assign po1603 = ~w6995;
assign po1604 = ~w6998;
assign po1605 = ~w7001;
assign po1606 = ~w7004;
assign po1607 = ~w7007;
assign po1608 = ~w7010;
assign po1609 = ~w7013;
assign po1610 = ~w7016;
assign po1611 = ~w7019;
assign po1612 = ~w7022;
assign po1613 = ~w7025;
assign po1614 = ~w7028;
assign po1615 = ~w7031;
assign po1616 = ~w7034;
assign po1617 = ~w7037;
assign po1618 = ~w7040;
assign po1619 = ~w7043;
assign po1620 = ~w7046;
assign po1621 = ~w7049;
assign po1622 = ~w7052;
assign po1623 = ~w7055;
assign po1624 = ~w7058;
assign po1625 = ~w7061;
assign po1626 = ~w7064;
assign po1627 = ~w7067;
assign po1628 = ~w7070;
assign po1629 = ~w7073;
assign po1630 = ~w7076;
assign po1631 = ~w7079;
assign po1632 = ~w7082;
assign po1633 = ~w7085;
assign po1634 = ~w7088;
assign po1635 = ~w7091;
assign po1636 = ~w7094;
assign po1637 = ~w7097;
assign po1638 = ~w7100;
assign po1639 = ~w7103;
assign po1640 = ~w7106;
assign po1641 = ~w7109;
assign po1642 = ~w7112;
assign po1643 = ~w7115;
assign po1644 = ~w7118;
assign po1645 = ~w7121;
assign po1646 = ~w7124;
assign po1647 = ~w7127;
assign po1648 = ~w7130;
assign po1649 = ~w7133;
assign po1650 = ~w7136;
assign po1651 = ~w7139;
assign po1652 = ~w7142;
assign po1653 = ~w7145;
assign po1654 = ~w7148;
assign po1655 = ~w7151;
assign po1656 = ~w7154;
assign po1657 = ~w7157;
assign po1658 = ~w7160;
assign po1659 = ~w7163;
assign po1660 = ~w7166;
assign po1661 = ~w7169;
assign po1662 = ~w7172;
assign po1663 = ~w7175;
assign po1664 = ~w7178;
assign po1665 = ~w7181;
assign po1666 = ~w7184;
assign po1667 = ~w7187;
assign po1668 = ~w7190;
assign po1669 = ~w7193;
assign po1670 = ~w7196;
assign po1671 = ~w7199;
assign po1672 = ~w7202;
assign po1673 = ~w7205;
assign po1674 = ~w7208;
assign po1675 = ~w7211;
assign po1676 = ~w7214;
assign po1677 = ~w7217;
assign po1678 = ~w7220;
assign po1679 = ~w7223;
assign po1680 = ~w7226;
assign po1681 = ~w7229;
assign po1682 = ~w7232;
assign po1683 = ~w7235;
assign po1684 = ~w7238;
assign po1685 = ~w7241;
assign po1686 = ~w7244;
assign po1687 = ~w7247;
assign po1688 = ~w7250;
assign po1689 = ~w7253;
assign po1690 = ~w7256;
assign po1691 = ~w7259;
assign po1692 = ~w7262;
assign po1693 = ~w7265;
assign po1694 = ~w7268;
assign po1695 = ~w7271;
assign po1696 = ~w7274;
assign po1697 = ~w7277;
assign po1698 = ~w7280;
assign po1699 = ~w7283;
assign po1700 = ~w7286;
assign po1701 = ~w7289;
assign po1702 = ~w7292;
assign po1703 = ~w7295;
assign po1704 = ~w7298;
assign po1705 = ~w7301;
assign po1706 = ~w7304;
assign po1707 = ~w7307;
assign po1708 = ~w7310;
assign po1709 = ~w7313;
assign po1710 = ~w7316;
assign po1711 = ~w7319;
assign po1712 = ~w7322;
assign po1713 = ~w7325;
assign po1714 = ~w7328;
assign po1715 = ~w7331;
assign po1716 = ~w7334;
assign po1717 = ~w7337;
assign po1718 = ~w7340;
assign po1719 = ~w7343;
assign po1720 = ~w7346;
assign po1721 = ~w7349;
assign po1722 = ~w7352;
assign po1723 = ~w7355;
assign po1724 = ~w7358;
assign po1725 = ~w7361;
assign po1726 = ~w7364;
assign po1727 = ~w7367;
assign po1728 = ~w7370;
assign po1729 = ~w7373;
assign po1730 = ~w7376;
assign po1731 = ~w7379;
assign po1732 = ~w7382;
assign po1733 = ~w7385;
assign po1734 = ~w7388;
assign po1735 = ~w7391;
assign po1736 = ~w7394;
assign po1737 = ~w7397;
assign po1738 = ~w7400;
assign po1739 = ~w7403;
assign po1740 = ~w7406;
assign po1741 = ~w7409;
assign po1742 = ~w7412;
assign po1743 = ~w7415;
assign po1744 = ~w7418;
assign po1745 = ~w7421;
assign po1746 = ~w7424;
assign po1747 = ~w7427;
assign po1748 = ~w7430;
assign po1749 = ~w7433;
assign po1750 = ~w7436;
assign po1751 = ~w7439;
assign po1752 = ~w7442;
assign po1753 = ~w7445;
assign po1754 = ~w7448;
assign po1755 = ~w7451;
assign po1756 = ~w7454;
assign po1757 = ~w7457;
assign po1758 = ~w7460;
assign po1759 = ~w7463;
assign po1760 = ~w7466;
assign po1761 = ~w7469;
assign po1762 = ~w7472;
assign po1763 = ~w7475;
assign po1764 = ~w7478;
assign po1765 = ~w7481;
assign po1766 = ~w7484;
assign po1767 = ~w7487;
assign po1768 = ~w7490;
assign po1769 = ~w7493;
assign po1770 = ~w7496;
assign po1771 = ~w7499;
assign po1772 = ~w7502;
assign po1773 = ~w7505;
assign po1774 = ~w7508;
assign po1775 = ~w7511;
assign po1776 = ~w7514;
assign po1777 = ~w7517;
assign po1778 = ~w7520;
assign po1779 = ~w7523;
assign po1780 = ~w7526;
assign po1781 = ~w7529;
assign po1782 = ~w7532;
assign po1783 = ~w7535;
assign po1784 = ~w7538;
assign po1785 = ~w7541;
assign po1786 = ~w7544;
assign po1787 = ~w7547;
assign po1788 = ~w7550;
assign po1789 = ~w7553;
assign po1790 = ~w7556;
assign po1791 = ~w7559;
assign po1792 = ~w7562;
assign po1793 = ~w7565;
assign po1794 = ~w7568;
assign po1795 = ~w7571;
assign po1796 = ~w7574;
assign po1797 = ~w7577;
assign po1798 = ~w7580;
assign po1799 = ~w7583;
assign po1800 = ~w7586;
assign po1801 = ~w7589;
assign po1802 = ~w7592;
assign po1803 = ~w7595;
assign po1804 = ~w7598;
assign po1805 = ~w7601;
assign po1806 = ~w7604;
assign po1807 = w7607;
assign po1808 = ~w7610;
assign po1809 = ~w7613;
assign po1810 = ~w7616;
assign po1811 = ~w7619;
assign po1812 = ~w7622;
assign po1813 = ~w7625;
assign po1814 = ~w7628;
assign po1815 = ~w7631;
assign po1816 = ~w7634;
assign po1817 = ~w7637;
assign po1818 = ~w7640;
assign po1819 = pi1880;
assign po1820 = ~w7643;
assign po1821 = ~w7646;
assign po1822 = ~w7649;
assign po1823 = ~w7652;
assign po1824 = ~w7655;
assign po1825 = ~w7658;
assign po1826 = ~w7661;
assign po1827 = ~w7664;
assign po1828 = ~w7667;
assign po1829 = ~w7670;
assign po1830 = ~w7673;
assign po1831 = ~w7676;
assign po1832 = ~w7679;
assign po1833 = ~w7682;
assign po1834 = ~w7685;
assign po1835 = ~w7688;
assign po1836 = ~w7691;
assign po1837 = ~w7694;
assign po1838 = ~w7697;
assign po1839 = ~w7700;
assign po1840 = ~w7703;
assign po1841 = ~w7706;
assign po1842 = ~w7709;
assign po1843 = ~w7712;
assign po1844 = ~w7715;
assign po1845 = ~w7718;
assign po1846 = ~w7721;
assign po1847 = ~w7724;
assign po1848 = ~w7727;
assign po1849 = ~w7730;
assign po1850 = ~w7733;
assign po1851 = ~w7736;
assign po1852 = ~w7739;
assign po1853 = ~w7742;
assign po1854 = ~w7745;
assign po1855 = ~w7748;
assign po1856 = ~w7751;
assign po1857 = ~w7754;
assign po1858 = ~w7757;
assign po1859 = ~w7760;
assign po1860 = ~w7763;
assign po1861 = ~w7766;
assign po1862 = ~w7769;
assign po1863 = ~w7772;
assign po1864 = ~w7775;
assign po1865 = ~w7778;
assign po1866 = ~w7781;
assign po1867 = ~w7784;
assign po1868 = ~w7787;
assign po1869 = ~w7790;
assign po1870 = ~w7793;
assign po1871 = ~w7796;
assign po1872 = ~w7799;
assign po1873 = ~w7802;
assign po1874 = ~w7805;
assign po1875 = ~w7808;
assign po1876 = ~w7811;
assign po1877 = ~w7814;
assign po1878 = ~w7817;
assign po1879 = ~w7820;
assign po1880 = ~w7823;
assign po1881 = ~w7826;
assign po1882 = ~w7829;
assign po1883 = ~w7833;
assign po1884 = ~w7836;
assign po1885 = w2400;
assign po1886 = ~w7854;
assign po1887 = ~w7871;
assign po1888 = ~w7888;
assign po1889 = ~w7891;
assign po1890 = ~w7894;
assign po1891 = ~w7897;
assign po1892 = ~w7900;
assign po1893 = ~w7903;
assign po1894 = ~w7906;
assign po1895 = ~w7909;
assign po1896 = ~w7912;
assign po1897 = ~w7915;
assign po1898 = ~w7918;
assign po1899 = ~w7921;
assign po1900 = ~w7924;
assign po1901 = ~w7927;
assign po1902 = ~w7930;
assign po1903 = ~w7933;
assign po1904 = ~w7936;
assign po1905 = ~w7939;
assign po1906 = ~w7942;
assign po1907 = ~w7945;
assign po1908 = ~w7948;
assign po1909 = ~w7965;
assign po1910 = ~w7982;
assign po1911 = ~w7999;
assign po1912 = ~w8016;
assign po1913 = ~w8033;
assign po1914 = ~w8050;
assign po1915 = ~w8067;
assign po1916 = ~w8084;
assign po1917 = ~w8101;
assign po1918 = ~w8118;
assign po1919 = ~w8135;
assign po1920 = ~w8152;
assign po1921 = ~w8155;
assign po1922 = ~w8158;
assign po1923 = ~w8161;
assign po1924 = ~w8164;
assign po1925 = ~w8167;
assign po1926 = ~w8170;
assign po1927 = w3365;
assign po1928 = ~w8173;
assign po1929 = w8175;
assign po1930 = w8176;
assign po1931 = pi1906;
assign po1932 = w3385;
assign po1933 = ~w8185;
assign po1934 = ~w8188;
assign po1935 = ~w8191;
assign po1936 = ~w8194;
assign po1937 = ~w8197;
assign po1938 = ~w8210;
assign po1939 = ~w8225;
assign po1940 = ~w8240;
assign po1941 = ~w8255;
assign po1942 = ~w8270;
assign po1943 = ~w8285;
assign po1944 = ~w8300;
assign po1945 = ~w8311;
assign po1946 = ~w8318;
assign po1947 = ~w8329;
assign po1948 = ~w8340;
assign po1949 = ~w8351;
assign po1950 = ~w8358;
assign po1951 = ~w8369;
assign po1952 = ~w8372;
assign po1953 = ~w8387;
assign po1954 = w8399;
assign po1955 = w8411;
assign po1956 = w5378;
assign po1957 = pi1928;
assign po1958 = w8423;
assign po1959 = w8434;
assign po1960 = w8446;
assign po1961 = w8458;
assign po1962 = w8464;
assign po1963 = w8470;
assign po1964 = ~w8472;
assign po1965 = ~w8474;
assign po1966 = w8478;
assign po1967 = w8484;
assign po1968 = w8488;
assign po1969 = w8491;
assign po1970 = w8494;
assign po1971 = w8498;
assign po1972 = w8501;
assign po1973 = ~w8504;
assign po1974 = ~w8507;
assign po1975 = ~w8510;
assign po1976 = ~w8513;
assign po1977 = ~w8516;
assign po1978 = ~w8518;
assign po1979 = pi1942;
assign po1980 = w8519;
assign po1981 = pi1953;
assign po1982 = pi1954;
assign po1983 = ~w8522;
assign po1984 = ~w8525;
assign po1985 = ~w8528;
assign po1986 = ~w8531;
assign po1987 = w8536;
assign po1988 = w8537;
assign po1989 = w8538;
assign po1990 = w8539;
assign po1991 = w8540;
assign po1992 = w8541;
assign po1993 = pi1992;
assign po1994 = pi1991;
assign po1995 = w8549;
assign po1996 = ~w8606;
assign po1997 = w8608;
assign po1998 = ~w8611;
assign po1999 = w8613;
assign po2000 = w8615;
assign po2001 = w8617;
assign po2002 = ~w8628;
assign po2003 = pi2011;
assign po2004 = pi2002;
assign po2005 = pi2012;
assign po2006 = w8637;
assign po2007 = w8644;
assign po2008 = w8647;
assign po2009 = ~w8650;
assign po2010 = ~w8653;
assign po2011 = ~w8656;
assign po2012 = ~w8659;
assign po2013 = ~w8662;
assign po2014 = w8664;
assign po2015 = w8666;
assign po2016 = w8668;
assign po2017 = w8670;
assign po2018 = w8672;
assign po2019 = w8674;
assign po2020 = w8676;
assign po2021 = w8678;
assign po2022 = w8680;
assign po2023 = w8682;
assign po2024 = w8684;
assign po2025 = w8686;
assign po2026 = w8688;
assign po2027 = w8690;
assign po2028 = w8692;
assign po2029 = ~w8695;
assign po2030 = ~w8698;
assign po2031 = ~w8701;
assign po2032 = ~w8704;
assign po2033 = w8706;
assign po2034 = ~w8709;
assign po2035 = ~w8712;
assign po2036 = ~w8716;
assign po2037 = w8719;
assign po2038 = ~w8721;
assign po2039 = ~w8723;
assign po2040 = w8724;
assign po2041 = w8727;
assign po2042 = pi2015;
assign po2043 = pi2014;
assign po2044 = ~w8730;
assign po2045 = ~w8734;
assign po2046 = w8736;
assign po2047 = w8739;
assign po2048 = ~w8742;
assign po2049 = ~w8745;
assign po2050 = ~w8746;
assign po2051 = ~w8749;
assign po2052 = w8752;
assign po2053 = ~w8758;
assign po2054 = w8761;
assign po2055 = ~w8763;
assign po2056 = ~w8765;
assign po2057 = ~w8767;
assign po2058 = ~w8769;
assign po2059 = w8776;
assign po2060 = w8788;
assign po2061 = w8800;
assign po2062 = pi2037;
assign po2063 = w8804;
assign po2064 = w8808;
assign po2065 = pi2081;
assign po2066 = w8812;
assign po2067 = w8815;
assign po2068 = w8818;
assign po2069 = w8826;
assign po2070 = w8827;
assign po2071 = w8828;
assign po2072 = ~w8838;
assign po2073 = ~w8845;
assign po2074 = ~w8852;
assign po2075 = ~w8859;
assign po2076 = ~w8866;
assign po2077 = ~w8873;
assign po2078 = ~w8880;
assign po2079 = ~w8887;
assign po2080 = ~w8894;
assign po2081 = ~w8901;
assign po2082 = w8902;
assign po2083 = w8906;
assign po2084 = w8907;
assign po2085 = w8908;
assign po2086 = w8913;
assign po2087 = w8914;
assign po2088 = ~w8917;
assign po2089 = ~w8924;
assign po2090 = ~w8931;
assign po2091 = ~w8938;
assign po2092 = ~w8945;
assign po2093 = ~w8952;
assign po2094 = ~w8959;
assign po2095 = ~w8966;
assign po2096 = ~w8973;
assign po2097 = ~w8980;
assign po2098 = ~w8987;
assign po2099 = ~w8994;
assign po2100 = ~w9001;
assign po2101 = ~w9008;
assign po2102 = ~w9015;
assign po2103 = ~w9022;
assign po2104 = ~w9029;
assign po2105 = ~w9036;
assign po2106 = w9037;
assign po2107 = w9041;
assign po2108 = w9043;
assign po2109 = w9047;
assign po2110 = w9049;
assign po2111 = w9051;
assign po2112 = ~w9061;
assign po2113 = ~w9068;
assign po2114 = ~w9075;
assign po2115 = ~w9082;
assign po2116 = ~w9089;
assign po2117 = ~w9096;
assign po2118 = ~w9103;
assign po2119 = ~w9110;
assign po2120 = ~w9117;
assign po2121 = ~w9124;
assign po2122 = ~w9131;
assign po2123 = ~w9138;
assign po2124 = ~w9145;
assign po2125 = ~w9152;
assign po2126 = ~w9159;
assign po2127 = ~w9166;
assign po2128 = ~w9173;
assign po2129 = ~w9180;
assign po2130 = ~w9187;
assign po2131 = ~w9194;
assign po2132 = pi2142;
assign po2133 = ~w9201;
assign po2134 = ~w9208;
assign po2135 = ~w9215;
assign po2136 = ~w9222;
assign po2137 = ~w9229;
assign po2138 = ~w9236;
assign po2139 = ~w9243;
assign po2140 = ~w9250;
assign po2141 = ~w9257;
assign po2142 = ~w9267;
assign po2143 = ~w9274;
assign po2144 = ~w9281;
assign po2145 = ~w9288;
assign po2146 = ~w9295;
assign po2147 = ~w9302;
assign po2148 = ~w9309;
assign po2149 = ~w9316;
assign po2150 = ~w9323;
assign po2151 = ~w9330;
assign po2152 = ~w9337;
assign po2153 = ~w9344;
assign po2154 = ~w9351;
assign po2155 = ~w9358;
assign po2156 = ~w9365;
assign po2157 = ~w9372;
assign po2158 = ~w9379;
assign po2159 = ~w9386;
assign po2160 = ~w9393;
assign po2161 = ~w9400;
assign po2162 = ~w9407;
assign po2163 = ~w9414;
assign po2164 = ~w9421;
assign po2165 = ~w9428;
assign po2166 = ~w9435;
assign po2167 = ~w9442;
assign po2168 = ~w9449;
assign po2169 = ~w9456;
assign po2170 = ~w9463;
assign po2171 = ~w9470;
assign po2172 = ~w9477;
assign po2173 = ~w9484;
assign po2174 = ~w9491;
assign po2175 = ~w9498;
assign po2176 = ~w9505;
assign po2177 = ~w9512;
assign po2178 = ~w9519;
assign po2179 = ~w9526;
assign po2180 = ~w9533;
assign po2181 = ~w9540;
assign po2182 = w684;
assign po2183 = w9541;
assign po2184 = ~w9544;
assign po2185 = w8634;
assign po2186 = w8782;
assign po2187 = w8794;
assign po2188 = w8823;
assign po2189 = w4989;
assign po2190 = w8417;
assign po2191 = w4963;
assign po2192 = w4976;
assign po2193 = pi2161;
assign po2194 = ~w9547;
assign po2195 = ~w9550;
assign po2196 = ~w9553;
assign po2197 = ~w9556;
assign po2198 = ~w9559;
assign po2199 = ~w9562;
assign po2200 = ~w9565;
assign po2201 = ~w9568;
assign po2202 = ~w9571;
assign po2203 = ~w9574;
assign po2204 = ~w9577;
assign po2205 = ~w9580;
assign po2206 = ~w9583;
assign po2207 = ~w9586;
assign po2208 = ~w9589;
assign po2209 = w9590;
assign po2210 = w5010;
assign po2211 = ~w9593;
assign po2212 = pi2164;
assign po2213 = w8533;
assign po2214 = ~pi2180;
assign po2215 = pi2165;
assign po2216 = ~pi2204;
assign po2217 = pi2205;
assign po2218 = pi2213;
assign po2219 = pi2210;
assign po2220 = pi2218;
assign po2221 = pi2230;
assign po2222 = pi2232;
assign po2223 = pi2229;
assign po2224 = pi2217;
assign po2225 = pi2237;
assign po2226 = pi2219;
assign po2227 = pi2235;
assign po2228 = pi2228;
assign po2229 = pi2236;
assign po2230 = pi2221;
assign po2231 = pi2225;
assign po2232 = pi2233;
assign po2233 = pi2234;
assign po2234 = pi2216;
assign po2235 = pi2212;
assign po2236 = pi2226;
assign po2237 = pi2206;
assign po2238 = pi2227;
assign po2239 = pi2211;
assign po2240 = pi2224;
assign po2241 = pi2231;
assign po2242 = pi2208;
assign po2243 = pi2215;
assign po2244 = pi2223;
assign po2245 = pi2209;
assign po2246 = pi2214;
assign po2247 = pi2222;
assign po2248 = pi2220;
assign po2249 = pi2207;
endmodule

module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970;
assign w0 = pi010 & pi013;
assign w1 = ~pi004 & ~pi006;
assign w2 = ~pi007 & ~pi008;
assign w3 = ~pi021 & w2;
assign w4 = w1 & w3;
assign w5 = w3 & w873;
assign w6 = pi007 & pi008;
assign w7 = ~pi010 & ~pi013;
assign w8 = w1 & w7;
assign w9 = ~pi014 & w8;
assign w10 = w8 & w874;
assign w11 = ~w5 & ~w10;
assign w12 = pi014 & ~w7;
assign w13 = ~pi016 & ~pi018;
assign w14 = ~pi017 & ~pi019;
assign w15 = ~pi009 & ~pi011;
assign w16 = ~pi005 & ~pi022;
assign w17 = w15 & w16;
assign w18 = w13 & w14;
assign w19 = w17 & w18;
assign w20 = (~pi012 & w2) | (~pi012 & w875) | (w2 & w875);
assign w21 = ~w12 & w20;
assign w22 = w19 & w21;
assign w23 = ~w11 & w22;
assign w24 = ~w15 & ~w16;
assign w25 = ~w17 & ~w24;
assign w26 = ~w23 & ~w25;
assign w27 = ~pi012 & ~pi014;
assign w28 = w3 & w27;
assign w29 = w8 & w19;
assign w30 = w28 & w29;
assign w31 = w29 & w876;
assign w32 = ~pi003 & ~pi129;
assign w33 = pi054 & w32;
assign w34 = (w33 & ~w25) | (w33 & w877) | (~w25 & w877);
assign w35 = ~w31 & w34;
assign w36 = ~w26 & w35;
assign w37 = ~pi054 & w32;
assign w38 = w32 & w878;
assign w39 = ~w36 & ~w38;
assign w40 = (w33 & ~w29) | (w33 & w879) | (~w29 & w879);
assign w41 = ~pi001 & w32;
assign w42 = ~w40 & ~w41;
assign w43 = ~pi011 & w27;
assign w44 = ~pi005 & ~pi009;
assign w45 = ~pi004 & w44;
assign w46 = w43 & w45;
assign w47 = ~pi006 & ~pi010;
assign w48 = ~w7 & ~w47;
assign w49 = w46 & ~w48;
assign w50 = pi012 & ~w44;
assign w51 = ~pi011 & ~w24;
assign w52 = ~w50 & w51;
assign w53 = w9 & w52;
assign w54 = ~w49 & ~w53;
assign w55 = (pi007 & ~w46) | (pi007 & w880) | (~w46 & w880);
assign w56 = ~pi021 & w14;
assign w57 = w14 & w881;
assign w58 = ~pi022 & w13;
assign w59 = w57 & w58;
assign w60 = ~w55 & w59;
assign w61 = ~pi001 & pi017;
assign w62 = pi054 & ~w61;
assign w63 = (w62 & ~w29) | (w62 & w882) | (~w29 & w882);
assign w64 = (w63 & w54) | (w63 & w883) | (w54 & w883);
assign w65 = ~w42 & ~w64;
assign w66 = ~pi046 & ~pi050;
assign w67 = ~pi043 & w66;
assign w68 = ~pi044 & ~pi045;
assign w69 = ~pi047 & ~pi048;
assign w70 = w68 & w69;
assign w71 = w67 & w70;
assign w72 = ~pi038 & ~pi040;
assign w73 = ~pi041 & ~pi042;
assign w74 = w72 & w73;
assign w75 = ~pi024 & ~pi049;
assign w76 = w74 & w75;
assign w77 = w71 & w76;
assign w78 = ~pi015 & ~pi020;
assign w79 = (pi082 & ~w77) | (pi082 & w884) | (~w77 & w884);
assign w80 = pi002 & w79;
assign w81 = ~pi049 & w71;
assign w82 = ~pi015 & ~pi024;
assign w83 = w74 & w82;
assign w84 = ~pi002 & ~pi020;
assign w85 = w74 & w885;
assign w86 = (pi082 & ~w81) | (pi082 & w886) | (~w81 & w886);
assign w87 = pi122 & pi127;
assign w88 = ~pi065 & ~w87;
assign w89 = pi002 & w87;
assign w90 = ~w88 & ~w89;
assign w91 = ~w86 & ~w90;
assign w92 = ~w80 & ~w91;
assign w93 = ~pi129 & ~w92;
assign w94 = pi000 & ~pi113;
assign w95 = ~pi123 & w94;
assign w96 = ~pi061 & ~pi118;
assign w97 = (w96 & ~w29) | (w96 & w887) | (~w29 & w887);
assign w98 = ~w95 & ~w97;
assign w99 = ~pi129 & ~w98;
assign w100 = ~pi013 & ~pi016;
assign w101 = w27 & w100;
assign w102 = w40 & w101;
assign w103 = ~pi004 & ~pi022;
assign w104 = w44 & w103;
assign w105 = ~pi011 & ~pi018;
assign w106 = w14 & w105;
assign w107 = w104 & w106;
assign w108 = w4 & w107;
assign w109 = w40 & w888;
assign w110 = w32 & w889;
assign w111 = ~w109 & ~w110;
assign w112 = w32 & w890;
assign w113 = w101 & w106;
assign w114 = w2 & w47;
assign w115 = w104 & w114;
assign w116 = w33 & w56;
assign w117 = w115 & w116;
assign w118 = ~pi029 & ~pi059;
assign w119 = ~pi025 & pi028;
assign w120 = w118 & w119;
assign w121 = w117 & w891;
assign w122 = ~w112 & ~w121;
assign w123 = w32 & w892;
assign w124 = pi025 & ~pi028;
assign w125 = w118 & w124;
assign w126 = w117 & w893;
assign w127 = ~w123 & ~w126;
assign w128 = w32 & w894;
assign w129 = w44 & w47;
assign w130 = w33 & ~w57;
assign w131 = ~pi021 & ~w6;
assign w132 = w103 & w131;
assign w133 = w129 & w132;
assign w134 = w133 & w895;
assign w135 = ~w128 & ~w134;
assign w136 = (~pi008 & ~w14) | (~pi008 & w896) | (~w14 & w896);
assign w137 = w27 & w938;
assign w138 = w13 & ~w56;
assign w139 = w115 & w138;
assign w140 = (pi054 & ~w139) | (pi054 & w897) | (~w139 & w897);
assign w141 = w32 & ~w136;
assign w142 = ~w140 & w141;
assign w143 = ~pi018 & w117;
assign w144 = w102 & w143;
assign w145 = w32 & w898;
assign w146 = ~w144 & ~w145;
assign w147 = w32 & w899;
assign w148 = w4 & w129;
assign w149 = w4 & w900;
assign w150 = ~pi011 & ~pi022;
assign w151 = ~pi012 & ~pi013;
assign w152 = ~pi017 & w151;
assign w153 = w13 & w150;
assign w154 = w152 & w153;
assign w155 = w149 & w154;
assign w156 = w40 & w155;
assign w157 = ~w147 & ~w156;
assign w158 = w32 & w901;
assign w159 = w113 & w148;
assign w160 = w40 & w159;
assign w161 = ~w158 & ~w160;
assign w162 = w32 & w902;
assign w163 = w43 & w117;
assign w164 = ~w30 & w163;
assign w165 = w100 & w164;
assign w166 = ~w162 & ~w165;
assign w167 = ~pi025 & ~pi028;
assign w168 = pi029 & ~pi059;
assign w169 = w167 & w168;
assign w170 = w117 & w903;
assign w171 = w32 & w904;
assign w172 = ~w170 & ~w171;
assign w173 = w32 & w905;
assign w174 = w13 & w164;
assign w175 = ~w173 & ~w174;
assign w176 = pi015 & w87;
assign w177 = ~pi070 & ~w87;
assign w178 = ~w176 & ~w177;
assign w179 = w81 & w83;
assign w180 = (pi082 & w77) | (pi082 & w906) | (w77 & w906);
assign w181 = ~w179 & w180;
assign w182 = (~pi129 & w86) | (~pi129 & w907) | (w86 & w907);
assign w183 = ~w181 & w182;
assign w184 = (pi016 & ~w32) | (pi016 & w908) | (~w32 & w908);
assign w185 = w15 & w103;
assign w186 = w56 & w185;
assign w187 = w101 & w114;
assign w188 = w186 & w187;
assign w189 = w7 & w33;
assign w190 = w28 & w189;
assign w191 = w107 & w190;
assign w192 = (~pi016 & ~w191) | (~pi016 & w909) | (~w191 & w909);
assign w193 = ~w184 & ~w192;
assign w194 = w32 & w910;
assign w195 = ~pi029 & pi059;
assign w196 = w167 & w195;
assign w197 = w117 & w911;
assign w198 = ~w194 & ~w197;
assign w199 = w32 & w912;
assign w200 = w137 & ~w188;
assign w201 = w143 & w200;
assign w202 = ~w199 & ~w201;
assign w203 = w32 & w913;
assign w204 = w58 & w137;
assign w205 = w130 & w204;
assign w206 = w149 & w205;
assign w207 = ~w203 & ~w206;
assign w208 = pi020 & w87;
assign w209 = ~pi071 & ~w87;
assign w210 = ~w208 & ~w209;
assign w211 = (pi020 & ~w81) | (pi020 & w914) | (~w81 & w914);
assign w212 = w79 & ~w211;
assign w213 = (~pi129 & w86) | (~pi129 & w915) | (w86 & w915);
assign w214 = ~w212 & w213;
assign w215 = w32 & w916;
assign w216 = ~pi014 & w154;
assign w217 = w130 & w216;
assign w218 = w148 & w217;
assign w219 = ~w215 & ~w218;
assign w220 = w32 & w917;
assign w221 = ~pi018 & w188;
assign w222 = w40 & w221;
assign w223 = ~w220 & ~w222;
assign w224 = ~pi023 & pi055;
assign w225 = pi061 & ~pi129;
assign w226 = ~w224 & w225;
assign w227 = pi024 & w87;
assign w228 = ~pi063 & ~w87;
assign w229 = ~w227 & ~w228;
assign w230 = w71 & w918;
assign w231 = (pi024 & ~w71) | (pi024 & w919) | (~w71 & w919);
assign w232 = pi082 & ~w230;
assign w233 = ~w231 & w232;
assign w234 = (~pi129 & w86) | (~pi129 & w920) | (w86 & w920);
assign w235 = ~w233 & w234;
assign w236 = ~pi053 & ~pi058;
assign w237 = ~pi085 & w236;
assign w238 = pi026 & ~pi027;
assign w239 = ~pi026 & pi027;
assign w240 = ~w238 & ~w239;
assign w241 = w237 & ~w240;
assign w242 = ~pi026 & ~pi027;
assign w243 = ~pi085 & w242;
assign w244 = ~pi053 & pi058;
assign w245 = w243 & w244;
assign w246 = ~w241 & ~w245;
assign w247 = pi053 & ~pi058;
assign w248 = w243 & w247;
assign w249 = w236 & w242;
assign w250 = pi085 & w249;
assign w251 = ~w248 & ~w250;
assign w252 = w246 & w251;
assign w253 = ~w252 & w921;
assign w254 = ~pi095 & ~pi100;
assign w255 = (~pi110 & ~w254) | (~pi110 & w922) | (~w254 & w922);
assign w256 = w237 & w242;
assign w257 = ~w255 & w256;
assign w258 = w256 & w923;
assign w259 = ~pi039 & ~pi051;
assign w260 = ~pi052 & w259;
assign w261 = w259 & w924;
assign w262 = w237 & w239;
assign w263 = w261 & w262;
assign w264 = w237 & w925;
assign w265 = ~w260 & w264;
assign w266 = ~pi085 & ~pi096;
assign w267 = ~pi110 & w266;
assign w268 = pi085 & pi116;
assign w269 = ~w267 & ~w268;
assign w270 = pi100 & w249;
assign w271 = ~w269 & w270;
assign w272 = ~w265 & ~w271;
assign w273 = ~w258 & ~w263;
assign w274 = w272 & w273;
assign w275 = ~w253 & w274;
assign w276 = w32 & ~w275;
assign w277 = ~w252 & w926;
assign w278 = w272 & ~w277;
assign w279 = w32 & ~w278;
assign w280 = ~w261 & w262;
assign w281 = ~pi100 & w249;
assign w282 = w249 & w927;
assign w283 = w266 & w928;
assign w284 = w281 & w283;
assign w285 = ~w280 & ~w282;
assign w286 = ~w284 & w285;
assign w287 = w32 & ~w286;
assign w288 = pi028 & ~pi116;
assign w289 = ~w282 & ~w288;
assign w290 = ~w252 & ~w289;
assign w291 = w256 & w929;
assign w292 = w260 & w264;
assign w293 = w262 & w930;
assign w294 = ~w284 & ~w291;
assign w295 = ~w292 & ~w293;
assign w296 = w294 & w295;
assign w297 = ~w290 & w296;
assign w298 = w32 & ~w297;
assign w299 = (~w257 & w252) | (~w257 & w931) | (w252 & w931);
assign w300 = pi029 & w32;
assign w301 = ~w299 & w300;
assign w302 = w243 & w932;
assign w303 = w266 & w933;
assign w304 = w281 & w303;
assign w305 = pi097 & w32;
assign w306 = (w305 & w304) | (w305 & w934) | (w304 & w934);
assign w307 = ~w301 & ~w306;
assign w308 = ~pi088 & pi106;
assign w309 = ~pi030 & ~pi109;
assign w310 = ~pi060 & pi109;
assign w311 = ~w309 & ~w310;
assign w312 = ~pi106 & ~w311;
assign w313 = ~pi129 & ~w308;
assign w314 = ~w312 & w313;
assign w315 = ~pi089 & pi106;
assign w316 = ~pi031 & ~pi109;
assign w317 = ~pi030 & pi109;
assign w318 = ~w316 & ~w317;
assign w319 = ~pi106 & ~w318;
assign w320 = ~pi129 & ~w315;
assign w321 = ~w319 & w320;
assign w322 = ~pi099 & pi106;
assign w323 = ~pi032 & ~pi109;
assign w324 = ~pi031 & pi109;
assign w325 = ~w323 & ~w324;
assign w326 = ~pi106 & ~w325;
assign w327 = ~pi129 & ~w322;
assign w328 = ~w326 & w327;
assign w329 = ~pi090 & pi106;
assign w330 = ~pi033 & ~pi109;
assign w331 = ~pi032 & pi109;
assign w332 = ~w330 & ~w331;
assign w333 = ~pi106 & ~w332;
assign w334 = ~pi129 & ~w329;
assign w335 = ~w333 & w334;
assign w336 = ~pi091 & pi106;
assign w337 = ~pi034 & ~pi109;
assign w338 = ~pi033 & pi109;
assign w339 = ~w337 & ~w338;
assign w340 = ~pi106 & ~w339;
assign w341 = ~pi129 & ~w336;
assign w342 = ~w340 & w341;
assign w343 = ~pi092 & pi106;
assign w344 = ~pi035 & ~pi109;
assign w345 = ~pi034 & pi109;
assign w346 = ~w344 & ~w345;
assign w347 = ~pi106 & ~w346;
assign w348 = ~pi129 & ~w343;
assign w349 = ~w347 & w348;
assign w350 = ~pi098 & pi106;
assign w351 = ~pi036 & ~pi109;
assign w352 = ~pi035 & pi109;
assign w353 = ~w351 & ~w352;
assign w354 = ~pi106 & ~w353;
assign w355 = ~pi129 & ~w350;
assign w356 = ~w354 & w355;
assign w357 = ~pi093 & pi106;
assign w358 = ~pi037 & ~pi109;
assign w359 = ~pi036 & pi109;
assign w360 = ~w358 & ~w359;
assign w361 = ~pi106 & ~w360;
assign w362 = ~pi129 & ~w357;
assign w363 = ~w361 & w362;
assign w364 = ~pi074 & ~w87;
assign w365 = pi038 & w87;
assign w366 = ~w364 & ~w365;
assign w367 = ~pi042 & ~pi044;
assign w368 = ~pi040 & w367;
assign w369 = (pi038 & ~w367) | (pi038 & w935) | (~w367 & w935);
assign w370 = w367 & w72;
assign w371 = ~w369 & ~w370;
assign w372 = w86 & w371;
assign w373 = (~pi129 & w86) | (~pi129 & w936) | (w86 & w936);
assign w374 = ~w372 & w373;
assign w375 = ~pi051 & pi109;
assign w376 = (pi039 & ~w375) | (pi039 & w937) | (~w375 & w937);
assign w377 = w259 & w939;
assign w378 = ~pi106 & ~w376;
assign w379 = ~w377 & w378;
assign w380 = ~pi129 & ~w379;
assign w381 = ~pi073 & ~w87;
assign w382 = pi040 & w87;
assign w383 = ~w381 & ~w382;
assign w384 = pi040 & ~w367;
assign w385 = ~w368 & ~w384;
assign w386 = w86 & w385;
assign w387 = (~pi129 & w86) | (~pi129 & w940) | (w86 & w940);
assign w388 = ~w386 & w387;
assign w389 = ~pi076 & ~w87;
assign w390 = pi041 & w87;
assign w391 = ~w389 & ~w390;
assign w392 = w66 & w370;
assign w393 = (pi041 & ~w370) | (pi041 & w941) | (~w370 & w941);
assign w394 = w370 & w942;
assign w395 = ~w393 & ~w394;
assign w396 = w86 & w395;
assign w397 = (~pi129 & w86) | (~pi129 & w943) | (w86 & w943);
assign w398 = ~w396 & w397;
assign w399 = ~pi072 & ~w87;
assign w400 = pi042 & w87;
assign w401 = ~w399 & ~w400;
assign w402 = pi042 & pi044;
assign w403 = ~w367 & ~w402;
assign w404 = w86 & w403;
assign w405 = (~pi129 & w86) | (~pi129 & w944) | (w86 & w944);
assign w406 = ~w404 & w405;
assign w407 = pi043 & ~w394;
assign w408 = w66 & w945;
assign w409 = w74 & w408;
assign w410 = pi082 & ~w409;
assign w411 = ~w407 & w410;
assign w412 = ~pi077 & ~w87;
assign w413 = pi043 & w87;
assign w414 = ~w412 & ~w413;
assign w415 = ~w86 & w414;
assign w416 = ~pi129 & ~w411;
assign w417 = ~w415 & w416;
assign w418 = ~pi067 & ~w87;
assign w419 = pi044 & w87;
assign w420 = ~w418 & ~w419;
assign w421 = ~w86 & w420;
assign w422 = (~pi129 & ~w86) | (~pi129 & w946) | (~w86 & w946);
assign w423 = ~w421 & w422;
assign w424 = ~pi047 & w409;
assign w425 = w409 & w69;
assign w426 = (pi045 & ~w409) | (pi045 & w947) | (~w409 & w947);
assign w427 = (pi082 & ~w71) | (pi082 & w948) | (~w71 & w948);
assign w428 = ~w426 & w427;
assign w429 = pi045 & w87;
assign w430 = ~pi068 & ~w87;
assign w431 = ~w429 & ~w430;
assign w432 = (~pi129 & w86) | (~pi129 & w949) | (w86 & w949);
assign w433 = ~w428 & w432;
assign w434 = pi046 & w87;
assign w435 = ~pi075 & ~w87;
assign w436 = ~w434 & ~w435;
assign w437 = ~pi050 & w370;
assign w438 = (pi046 & ~w370) | (pi046 & w950) | (~w370 & w950);
assign w439 = ~w392 & ~w438;
assign w440 = w86 & w439;
assign w441 = (~pi129 & w86) | (~pi129 & w951) | (w86 & w951);
assign w442 = ~w440 & w441;
assign w443 = ~pi064 & ~w87;
assign w444 = pi047 & w87;
assign w445 = ~w443 & ~w444;
assign w446 = pi047 & ~w409;
assign w447 = ~w424 & ~w446;
assign w448 = w86 & w447;
assign w449 = (~pi129 & w86) | (~pi129 & w952) | (w86 & w952);
assign w450 = ~w448 & w449;
assign w451 = pi048 & w87;
assign w452 = ~pi062 & ~w87;
assign w453 = ~w451 & ~w452;
assign w454 = ~w86 & w453;
assign w455 = (pi048 & ~w409) | (pi048 & w953) | (~w409 & w953);
assign w456 = w86 & w954;
assign w457 = ~pi129 & ~w454;
assign w458 = ~w456 & w457;
assign w459 = pi049 & w87;
assign w460 = ~pi069 & ~w87;
assign w461 = ~w459 & ~w460;
assign w462 = pi049 & ~w230;
assign w463 = ~w77 & w86;
assign w464 = ~w462 & w463;
assign w465 = (~pi129 & w86) | (~pi129 & w955) | (w86 & w955);
assign w466 = ~w464 & w465;
assign w467 = ~pi066 & ~w87;
assign w468 = pi050 & w87;
assign w469 = ~w467 & ~w468;
assign w470 = pi050 & ~w370;
assign w471 = ~w437 & ~w470;
assign w472 = w86 & w471;
assign w473 = (~pi129 & w86) | (~pi129 & w956) | (w86 & w956);
assign w474 = ~w472 & w473;
assign w475 = pi051 & ~pi109;
assign w476 = ~pi106 & ~w375;
assign w477 = ~w475 & w476;
assign w478 = ~pi129 & ~w477;
assign w479 = pi052 & ~w375;
assign w480 = (~pi106 & ~w375) | (~pi106 & w957) | (~w375 & w957);
assign w481 = ~w479 & w480;
assign w482 = ~pi129 & ~w481;
assign w483 = ~pi116 & w32;
assign w484 = w248 & w483;
assign w485 = ~w306 & ~w484;
assign w486 = ~w86 & ~w87;
assign w487 = ~pi129 & ~w486;
assign w488 = ~pi123 & ~pi129;
assign w489 = pi114 & ~pi122;
assign w490 = w488 & w489;
assign w491 = ~w245 & ~w264;
assign w492 = pi094 & ~w491;
assign w493 = pi037 & ~pi116;
assign w494 = w237 & w958;
assign w495 = ~w241 & ~w249;
assign w496 = ~pi026 & pi037;
assign w497 = (w496 & ~w495) | (w496 & w959) | (~w495 & w959);
assign w498 = ~w302 & ~w494;
assign w499 = ~w492 & w498;
assign w500 = ~w497 & w499;
assign w501 = w32 & ~w500;
assign w502 = w243 & w960;
assign w503 = w495 & w961;
assign w504 = pi060 & w302;
assign w505 = (~w504 & w503) | (~w504 & w962) | (w503 & w962);
assign w506 = w32 & ~w505;
assign w507 = pi058 & ~pi116;
assign w508 = (~w507 & ~w262) | (~w507 & w963) | (~w262 & w963);
assign w509 = ~w292 & w508;
assign w510 = w32 & ~w246;
assign w511 = ~w509 & w510;
assign w512 = pi059 & w32;
assign w513 = ~w299 & w512;
assign w514 = w32 & w255;
assign w515 = w256 & w514;
assign w516 = pi096 & w515;
assign w517 = ~w513 & ~w516;
assign w518 = ~pi117 & ~pi122;
assign w519 = pi123 & w518;
assign w520 = pi060 & ~w518;
assign w521 = ~w519 & ~w520;
assign w522 = ~pi114 & ~pi122;
assign w523 = pi123 & ~pi129;
assign w524 = w522 & w523;
assign w525 = pi131 & pi132;
assign w526 = pi133 & w525;
assign w527 = w525 & w964;
assign w528 = ~pi137 & ~pi138;
assign w529 = pi140 & w528;
assign w530 = w527 & w529;
assign w531 = w527 & w528;
assign w532 = (~pi062 & ~w527) | (~pi062 & w965) | (~w527 & w965);
assign w533 = ~pi129 & ~w530;
assign w534 = ~w532 & w533;
assign w535 = pi142 & w528;
assign w536 = w527 & w535;
assign w537 = (~pi063 & ~w527) | (~pi063 & w966) | (~w527 & w966);
assign w538 = ~pi129 & ~w536;
assign w539 = ~w537 & w538;
assign w540 = pi139 & w528;
assign w541 = w527 & w540;
assign w542 = (~pi064 & ~w527) | (~pi064 & w967) | (~w527 & w967);
assign w543 = ~pi129 & ~w541;
assign w544 = ~w542 & w543;
assign w545 = pi146 & w528;
assign w546 = w527 & w545;
assign w547 = (~pi065 & ~w527) | (~pi065 & w968) | (~w527 & w968);
assign w548 = ~pi129 & ~w546;
assign w549 = ~w547 & w548;
assign w550 = w525 & w969;
assign w551 = pi143 & w528;
assign w552 = w550 & w551;
assign w553 = w528 & w550;
assign w554 = (~pi066 & ~w550) | (~pi066 & w970) | (~w550 & w970);
assign w555 = ~pi129 & ~w552;
assign w556 = ~w554 & w555;
assign w557 = w540 & w550;
assign w558 = ~pi067 & ~w553;
assign w559 = ~pi129 & ~w557;
assign w560 = ~w558 & w559;
assign w561 = pi141 & w528;
assign w562 = w527 & w561;
assign w563 = ~pi068 & ~w531;
assign w564 = ~pi129 & ~w562;
assign w565 = ~w563 & w564;
assign w566 = w527 & w551;
assign w567 = ~pi069 & ~w531;
assign w568 = ~pi129 & ~w566;
assign w569 = ~w567 & w568;
assign w570 = pi144 & w528;
assign w571 = w527 & w570;
assign w572 = ~pi070 & ~w531;
assign w573 = ~pi129 & ~w571;
assign w574 = ~w572 & w573;
assign w575 = pi145 & w528;
assign w576 = w527 & w575;
assign w577 = ~pi071 & ~w531;
assign w578 = ~pi129 & ~w576;
assign w579 = ~w577 & w578;
assign w580 = w529 & w550;
assign w581 = ~pi072 & ~w553;
assign w582 = ~pi129 & ~w580;
assign w583 = ~w581 & w582;
assign w584 = w550 & w561;
assign w585 = ~pi073 & ~w553;
assign w586 = ~pi129 & ~w584;
assign w587 = ~w585 & w586;
assign w588 = w535 & w550;
assign w589 = ~pi074 & ~w553;
assign w590 = ~pi129 & ~w588;
assign w591 = ~w589 & w590;
assign w592 = w550 & w570;
assign w593 = ~pi075 & ~w553;
assign w594 = ~pi129 & ~w592;
assign w595 = ~w593 & w594;
assign w596 = w550 & w575;
assign w597 = ~pi076 & ~w553;
assign w598 = ~pi129 & ~w596;
assign w599 = ~w597 & w598;
assign w600 = w545 & w550;
assign w601 = ~pi077 & ~w553;
assign w602 = ~pi129 & ~w600;
assign w603 = ~w601 & w602;
assign w604 = pi137 & ~pi138;
assign w605 = ~pi142 & w604;
assign w606 = w550 & w605;
assign w607 = w550 & w604;
assign w608 = ~pi078 & ~w607;
assign w609 = ~pi129 & ~w606;
assign w610 = ~w608 & w609;
assign w611 = ~pi143 & w604;
assign w612 = w550 & w611;
assign w613 = ~pi079 & ~w607;
assign w614 = ~pi129 & ~w612;
assign w615 = ~w613 & w614;
assign w616 = ~pi144 & w604;
assign w617 = w550 & w616;
assign w618 = ~pi080 & ~w607;
assign w619 = ~pi129 & ~w617;
assign w620 = ~w618 & w619;
assign w621 = ~pi145 & w604;
assign w622 = w550 & w621;
assign w623 = ~pi081 & ~w607;
assign w624 = ~pi129 & ~w622;
assign w625 = ~w623 & w624;
assign w626 = ~pi146 & w604;
assign w627 = w550 & w626;
assign w628 = ~pi082 & ~w607;
assign w629 = ~pi129 & ~w627;
assign w630 = ~w628 & w629;
assign w631 = ~pi137 & pi138;
assign w632 = pi089 & w631;
assign w633 = pi031 & w604;
assign w634 = ~pi062 & w528;
assign w635 = ~w632 & ~w633;
assign w636 = ~w634 & w635;
assign w637 = pi136 & ~w636;
assign w638 = ~pi136 & w631;
assign w639 = pi119 & w638;
assign w640 = pi072 & ~pi137;
assign w641 = ~pi136 & ~w631;
assign w642 = pi115 & pi138;
assign w643 = ~pi087 & w604;
assign w644 = ~w640 & ~w642;
assign w645 = w641 & w644;
assign w646 = ~w643 & w645;
assign w647 = ~w639 & ~w646;
assign w648 = ~w637 & w647;
assign w649 = ~pi141 & w604;
assign w650 = w550 & w649;
assign w651 = ~pi084 & ~w607;
assign w652 = ~pi129 & ~w650;
assign w653 = ~w651 & w652;
assign w654 = w250 & w483;
assign w655 = ~w516 & ~w654;
assign w656 = ~pi139 & w604;
assign w657 = w550 & w656;
assign w658 = ~pi086 & ~w607;
assign w659 = ~pi129 & ~w657;
assign w660 = ~w658 & w659;
assign w661 = ~pi140 & w604;
assign w662 = w550 & w661;
assign w663 = ~pi087 & ~w607;
assign w664 = ~pi129 & ~w662;
assign w665 = ~w663 & w664;
assign w666 = w527 & w656;
assign w667 = w527 & w604;
assign w668 = ~pi088 & ~w667;
assign w669 = ~pi129 & ~w666;
assign w670 = ~w668 & w669;
assign w671 = w527 & w661;
assign w672 = ~pi089 & ~w667;
assign w673 = ~pi129 & ~w671;
assign w674 = ~w672 & w673;
assign w675 = w527 & w605;
assign w676 = ~pi090 & ~w667;
assign w677 = ~pi129 & ~w675;
assign w678 = ~w676 & w677;
assign w679 = w527 & w611;
assign w680 = ~pi091 & ~w667;
assign w681 = ~pi129 & ~w679;
assign w682 = ~w680 & w681;
assign w683 = w527 & w616;
assign w684 = ~pi092 & ~w667;
assign w685 = ~pi129 & ~w683;
assign w686 = ~w684 & w685;
assign w687 = w527 & w626;
assign w688 = ~pi093 & ~w667;
assign w689 = ~pi129 & ~w687;
assign w690 = ~w688 & w689;
assign w691 = pi082 & w638;
assign w692 = w526 & w691;
assign w693 = ~pi094 & ~w692;
assign w694 = ~pi142 & w692;
assign w695 = ~pi129 & ~w693;
assign w696 = ~w694 & w695;
assign w697 = ~pi003 & ~pi110;
assign w698 = ~w526 & ~w697;
assign w699 = ~w692 & ~w698;
assign w700 = pi095 & w699;
assign w701 = pi143 & w692;
assign w702 = ~w700 & ~w701;
assign w703 = ~pi129 & ~w702;
assign w704 = pi096 & w699;
assign w705 = pi146 & w692;
assign w706 = ~w704 & ~w705;
assign w707 = ~pi129 & ~w706;
assign w708 = pi097 & w699;
assign w709 = pi145 & w692;
assign w710 = ~w708 & ~w709;
assign w711 = ~pi129 & ~w710;
assign w712 = w527 & w621;
assign w713 = ~pi098 & ~w667;
assign w714 = ~pi129 & ~w712;
assign w715 = ~w713 & w714;
assign w716 = w527 & w649;
assign w717 = ~pi099 & ~w667;
assign w718 = ~pi129 & ~w716;
assign w719 = ~w717 & w718;
assign w720 = pi100 & w699;
assign w721 = pi144 & w692;
assign w722 = ~w720 & ~w721;
assign w723 = ~pi129 & ~w722;
assign w724 = pi137 & pi138;
assign w725 = pi096 & w724;
assign w726 = pi082 & w604;
assign w727 = ~pi077 & w528;
assign w728 = pi124 & w631;
assign w729 = ~pi136 & ~w725;
assign w730 = ~w726 & ~w727;
assign w731 = ~w728 & w730;
assign w732 = w729 & w731;
assign w733 = pi093 & w631;
assign w734 = ~pi065 & w528;
assign w735 = pi037 & w604;
assign w736 = pi136 & ~w733;
assign w737 = ~w734 & ~w735;
assign w738 = w736 & w737;
assign w739 = ~w732 & ~w738;
assign w740 = pi091 & w631;
assign w741 = ~pi069 & w528;
assign w742 = pi034 & w604;
assign w743 = ~w740 & ~w741;
assign w744 = ~w742 & w743;
assign w745 = pi136 & ~w744;
assign w746 = ~pi079 & w604;
assign w747 = ~pi066 & ~pi138;
assign w748 = ~pi095 & pi138;
assign w749 = pi137 & ~w748;
assign w750 = ~w747 & ~w749;
assign w751 = ~pi136 & ~w746;
assign w752 = ~w750 & w751;
assign w753 = ~w745 & ~w752;
assign w754 = pi090 & w631;
assign w755 = ~pi063 & w528;
assign w756 = pi033 & w604;
assign w757 = ~w754 & ~w755;
assign w758 = ~w756 & w757;
assign w759 = pi136 & ~w758;
assign w760 = ~pi094 & pi138;
assign w761 = ~pi078 & w604;
assign w762 = pi074 & ~pi137;
assign w763 = ~w760 & ~w762;
assign w764 = w641 & w763;
assign w765 = ~w761 & w764;
assign w766 = ~w759 & ~w765;
assign w767 = pi032 & w604;
assign w768 = ~pi068 & w528;
assign w769 = pi099 & w631;
assign w770 = ~w767 & ~w768;
assign w771 = ~w769 & w770;
assign w772 = pi136 & ~w771;
assign w773 = pi073 & ~pi137;
assign w774 = ~pi084 & w604;
assign w775 = pi112 & pi138;
assign w776 = ~w773 & ~w775;
assign w777 = w641 & w776;
assign w778 = ~w774 & w777;
assign w779 = ~w772 & ~w778;
assign w780 = pi125 & w631;
assign w781 = pi080 & w604;
assign w782 = ~pi075 & w528;
assign w783 = pi100 & w724;
assign w784 = ~pi136 & ~w780;
assign w785 = ~w781 & ~w782;
assign w786 = ~w783 & w785;
assign w787 = w784 & w786;
assign w788 = ~pi070 & w528;
assign w789 = pi035 & w604;
assign w790 = pi092 & w631;
assign w791 = pi136 & ~w788;
assign w792 = ~w789 & ~w790;
assign w793 = w791 & w792;
assign w794 = ~w787 & ~w793;
assign w795 = pi116 & w32;
assign w796 = pi085 & w795;
assign w797 = ~w515 & ~w796;
assign w798 = ~pi071 & w528;
assign w799 = pi036 & w604;
assign w800 = pi098 & w631;
assign w801 = ~w798 & ~w799;
assign w802 = ~w800 & w801;
assign w803 = pi136 & ~w802;
assign w804 = ~pi023 & w631;
assign w805 = ~pi097 & w724;
assign w806 = ~pi081 & w604;
assign w807 = pi076 & w528;
assign w808 = ~pi136 & ~w804;
assign w809 = ~w805 & ~w806;
assign w810 = ~w807 & w809;
assign w811 = w808 & w810;
assign w812 = ~w803 & ~w811;
assign w813 = ~pi064 & w528;
assign w814 = pi030 & w604;
assign w815 = pi088 & w631;
assign w816 = ~w813 & ~w814;
assign w817 = ~w815 & w816;
assign w818 = pi136 & ~w817;
assign w819 = ~pi120 & w631;
assign w820 = ~pi111 & w724;
assign w821 = pi067 & w528;
assign w822 = ~pi086 & w604;
assign w823 = ~pi136 & ~w819;
assign w824 = ~w820 & ~w821;
assign w825 = ~w822 & w824;
assign w826 = w823 & w825;
assign w827 = ~w818 & ~w826;
assign w828 = ~pi026 & w260;
assign w829 = ~w240 & w795;
assign w830 = ~w828 & w829;
assign w831 = ~pi097 & w244;
assign w832 = ~w247 & ~w831;
assign w833 = w795 & ~w832;
assign w834 = ~pi129 & w526;
assign w835 = ~pi111 & ~w691;
assign w836 = ~pi139 & w691;
assign w837 = w834 & ~w835;
assign w838 = ~w836 & w837;
assign w839 = ~pi141 & w691;
assign w840 = pi112 & ~w691;
assign w841 = w834 & ~w839;
assign w842 = ~w840 & w841;
assign w843 = w33 & ~w150;
assign w844 = ~pi113 & w37;
assign w845 = ~w843 & ~w844;
assign w846 = ~pi140 & w691;
assign w847 = pi115 & ~w691;
assign w848 = w834 & ~w846;
assign w849 = ~w847 & w848;
assign w850 = ~pi004 & ~pi007;
assign w851 = ~pi009 & ~pi012;
assign w852 = w850 & w851;
assign w853 = w33 & ~w852;
assign w854 = pi122 & ~pi129;
assign w855 = ~pi054 & ~pi118;
assign w856 = pi054 & ~w169;
assign w857 = ~pi129 & ~w855;
assign w858 = ~w856 & w857;
assign w859 = ~pi129 & ~w254;
assign w860 = ~pi120 & w697;
assign w861 = ~pi111 & ~pi129;
assign w862 = ~w860 & w861;
assign w863 = pi081 & pi120;
assign w864 = ~pi129 & w863;
assign w865 = ~pi129 & ~pi134;
assign w866 = ~pi129 & ~pi135;
assign w867 = pi057 & ~pi129;
assign w868 = ~pi096 & pi125;
assign w869 = ~pi003 & ~w868;
assign w870 = ~pi129 & ~w869;
assign w871 = ~pi126 & pi132;
assign w872 = pi133 & w871;
assign w873 = w1 & ~w0;
assign w874 = ~pi014 & ~w6;
assign w875 = ~pi021 & ~pi012;
assign w876 = w28 & pi000;
assign w877 = ~pi056 & w33;
assign w878 = ~pi054 & ~pi000;
assign w879 = ~w28 & w33;
assign w880 = ~w8 & pi007;
assign w881 = ~pi021 & ~pi008;
assign w882 = ~w28 & w62;
assign w883 = ~w60 & w63;
assign w884 = ~w78 & pi082;
assign w885 = w82 & w84;
assign w886 = ~w85 & pi082;
assign w887 = ~w28 & w96;
assign w888 = w101 & w108;
assign w889 = ~pi054 & pi004;
assign w890 = ~pi054 & pi005;
assign w891 = w113 & w120;
assign w892 = ~pi054 & pi006;
assign w893 = w113 & w125;
assign w894 = ~pi054 & pi007;
assign w895 = w113 & w130;
assign w896 = ~pi054 & ~pi008;
assign w897 = ~w137 & pi054;
assign w898 = ~pi054 & pi009;
assign w899 = ~pi054 & pi010;
assign w900 = w129 & ~pi019;
assign w901 = ~pi054 & pi011;
assign w902 = ~pi054 & pi012;
assign w903 = w113 & w169;
assign w904 = ~pi054 & pi013;
assign w905 = ~pi054 & pi014;
assign w906 = ~pi015 & pi082;
assign w907 = ~w178 & ~pi129;
assign w908 = pi054 & pi016;
assign w909 = w188 & ~pi016;
assign w910 = ~pi054 & pi017;
assign w911 = w113 & w196;
assign w912 = ~pi054 & pi018;
assign w913 = ~pi054 & pi019;
assign w914 = ~w83 & pi020;
assign w915 = ~w210 & ~pi129;
assign w916 = ~pi054 & pi021;
assign w917 = ~pi054 & pi022;
assign w918 = w74 & ~pi024;
assign w919 = ~w74 & pi024;
assign w920 = ~w229 & ~pi129;
assign w921 = ~pi116 & pi025;
assign w922 = pi097 & ~pi110;
assign w923 = ~w255 & pi025;
assign w924 = ~pi052 & pi116;
assign w925 = w238 & pi116;
assign w926 = ~pi116 & pi026;
assign w927 = ~pi100 & w268;
assign w928 = ~pi110 & pi095;
assign w929 = ~w255 & pi028;
assign w930 = ~w261 & pi116;
assign w931 = pi116 & ~w257;
assign w932 = w244 & pi116;
assign w933 = ~pi110 & ~pi095;
assign w934 = w302 & w305;
assign w935 = pi040 & pi038;
assign w936 = ~w366 & ~pi129;
assign w937 = pi052 & pi039;
assign w938 = ~pi011 & ~pi013;
assign w939 = ~pi052 & pi109;
assign w940 = ~w383 & ~pi129;
assign w941 = ~w66 & pi041;
assign w942 = w66 & ~pi041;
assign w943 = ~w391 & ~pi129;
assign w944 = ~w401 & ~pi129;
assign w945 = ~pi043 & ~pi044;
assign w946 = ~pi044 & ~pi129;
assign w947 = ~w69 & pi045;
assign w948 = ~w74 & pi082;
assign w949 = ~w431 & ~pi129;
assign w950 = pi050 & pi046;
assign w951 = ~w436 & ~pi129;
assign w952 = ~w445 & ~pi129;
assign w953 = pi047 & pi048;
assign w954 = ~w425 & ~w455;
assign w955 = ~w461 & ~pi129;
assign w956 = ~w469 & ~pi129;
assign w957 = pi052 & ~pi106;
assign w958 = w238 & w493;
assign w959 = w248 & w496;
assign w960 = w244 & ~pi116;
assign w961 = ~w248 & ~w502;
assign w962 = ~pi057 & ~w504;
assign w963 = ~w261 & ~w507;
assign w964 = pi133 & pi136;
assign w965 = ~w528 & ~pi062;
assign w966 = ~w528 & ~pi063;
assign w967 = ~w528 & ~pi064;
assign w968 = ~w528 & ~pi065;
assign w969 = pi133 & ~pi136;
assign w970 = ~w528 & ~pi066;
assign one = 1;
assign po000 = pi108;
assign po001 = pi083;
assign po002 = pi104;
assign po003 = pi103;
assign po004 = pi102;
assign po005 = pi105;
assign po006 = pi107;
assign po007 = pi101;
assign po008 = pi126;
assign po009 = pi121;
assign po010 = pi001;
assign po011 = pi000;
assign po012 = one;
assign po013 = pi130;
assign po014 = pi128;
assign po015 = w39;
assign po016 = ~w65;
assign po017 = w93;
assign po018 = w99;
assign po019 = ~w111;
assign po020 = ~w122;
assign po021 = ~w127;
assign po022 = ~w135;
assign po023 = w142;
assign po024 = ~w146;
assign po025 = ~w157;
assign po026 = ~w161;
assign po027 = ~w166;
assign po028 = ~w172;
assign po029 = ~w175;
assign po030 = w183;
assign po031 = w193;
assign po032 = ~w198;
assign po033 = ~w202;
assign po034 = ~w207;
assign po035 = w214;
assign po036 = ~w219;
assign po037 = ~w223;
assign po038 = w226;
assign po039 = w235;
assign po040 = w276;
assign po041 = w279;
assign po042 = w287;
assign po043 = w298;
assign po044 = ~w307;
assign po045 = w314;
assign po046 = w321;
assign po047 = w328;
assign po048 = w335;
assign po049 = w342;
assign po050 = w349;
assign po051 = w356;
assign po052 = w363;
assign po053 = w374;
assign po054 = w380;
assign po055 = w388;
assign po056 = w398;
assign po057 = w406;
assign po058 = w417;
assign po059 = w423;
assign po060 = w433;
assign po061 = w442;
assign po062 = w450;
assign po063 = w458;
assign po064 = w466;
assign po065 = w474;
assign po066 = w478;
assign po067 = w482;
assign po068 = ~w485;
assign po069 = ~w487;
assign po070 = w490;
assign po071 = w501;
assign po072 = w506;
assign po073 = w511;
assign po074 = ~w517;
assign po075 = ~w521;
assign po076 = w524;
assign po077 = ~w534;
assign po078 = ~w539;
assign po079 = ~w544;
assign po080 = ~w549;
assign po081 = ~w556;
assign po082 = ~w560;
assign po083 = ~w565;
assign po084 = ~w569;
assign po085 = ~w574;
assign po086 = ~w579;
assign po087 = ~w583;
assign po088 = ~w587;
assign po089 = ~w591;
assign po090 = ~w595;
assign po091 = ~w599;
assign po092 = ~w603;
assign po093 = w610;
assign po094 = w615;
assign po095 = w620;
assign po096 = w625;
assign po097 = w630;
assign po098 = ~w648;
assign po099 = w653;
assign po100 = ~w655;
assign po101 = w660;
assign po102 = w665;
assign po103 = w670;
assign po104 = w674;
assign po105 = w678;
assign po106 = w682;
assign po107 = w686;
assign po108 = w690;
assign po109 = w696;
assign po110 = w703;
assign po111 = w707;
assign po112 = w711;
assign po113 = w715;
assign po114 = w719;
assign po115 = w723;
assign po116 = w739;
assign po117 = ~w753;
assign po118 = ~w766;
assign po119 = ~w779;
assign po120 = w794;
assign po121 = ~w797;
assign po122 = ~w812;
assign po123 = ~w827;
assign po124 = w830;
assign po125 = w833;
assign po126 = w838;
assign po127 = w842;
assign po128 = ~w845;
assign po129 = ~w488;
assign po130 = w849;
assign po131 = w853;
assign po132 = ~w854;
assign po133 = w858;
assign po134 = w859;
assign po135 = w862;
assign po136 = w864;
assign po137 = ~w865;
assign po138 = ~w866;
assign po139 = w867;
assign po140 = w870;
assign po141 = w872;
endmodule

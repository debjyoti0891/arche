module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492;
assign w0 = pi046 & ~pi054;
assign w1 = pi045 & ~pi053;
assign w2 = ~w0 & ~w1;
assign w3 = ~pi045 & pi053;
assign w4 = ~pi044 & pi052;
assign w5 = ~w3 & ~w4;
assign w6 = ~w2 & w5;
assign w7 = pi044 & ~pi052;
assign w8 = pi043 & ~pi051;
assign w9 = ~w7 & ~w8;
assign w10 = ~w6 & w9;
assign w11 = ~pi042 & pi050;
assign w12 = ~pi041 & pi049;
assign w13 = ~pi040 & pi048;
assign w14 = ~w12 & ~w13;
assign w15 = ~pi043 & pi051;
assign w16 = ~w11 & ~w15;
assign w17 = w14 & w16;
assign w18 = ~w10 & w17;
assign w19 = pi039 & ~pi047;
assign w20 = pi042 & ~pi050;
assign w21 = pi041 & ~pi049;
assign w22 = ~w20 & ~w21;
assign w23 = w14 & ~w22;
assign w24 = pi040 & ~pi048;
assign w25 = ~w19 & ~w24;
assign w26 = ~w23 & w25;
assign w27 = ~w18 & w26;
assign w28 = ~pi039 & pi047;
assign w29 = ~w27 & ~w28;
assign w30 = pi002 & w29;
assign w31 = pi040 & ~pi216;
assign w32 = pi039 & ~pi215;
assign w33 = ~w31 & ~w32;
assign w34 = ~pi039 & pi215;
assign w35 = ~w33 & ~w34;
assign w36 = ~pi043 & pi219;
assign w37 = ~pi042 & pi218;
assign w38 = ~w36 & ~w37;
assign w39 = pi042 & ~pi218;
assign w40 = pi041 & ~pi217;
assign w41 = ~w39 & ~w40;
assign w42 = ~w38 & w41;
assign w43 = pi046 & ~pi222;
assign w44 = pi045 & ~pi221;
assign w45 = ~w43 & ~w44;
assign w46 = ~pi045 & pi221;
assign w47 = ~pi044 & pi220;
assign w48 = ~w46 & ~w47;
assign w49 = ~w45 & w48;
assign w50 = pi044 & ~pi220;
assign w51 = pi043 & ~pi219;
assign w52 = ~w50 & ~w51;
assign w53 = w41 & w52;
assign w54 = ~w49 & w53;
assign w55 = ~w42 & ~w54;
assign w56 = ~pi041 & pi217;
assign w57 = ~pi040 & pi216;
assign w58 = ~w56 & ~w57;
assign w59 = ~w34 & w58;
assign w60 = ~w54 & w16168;
assign w61 = ~w35 & ~w60;
assign w62 = pi039 & ~pi223;
assign w63 = ~pi045 & pi229;
assign w64 = pi046 & ~pi230;
assign w65 = ~w63 & w64;
assign w66 = pi045 & ~pi229;
assign w67 = pi044 & ~pi228;
assign w68 = ~w66 & ~w67;
assign w69 = ~w65 & w68;
assign w70 = ~pi042 & pi226;
assign w71 = ~pi044 & pi228;
assign w72 = ~pi043 & pi227;
assign w73 = ~w70 & ~w71;
assign w74 = ~w72 & w73;
assign w75 = ~w69 & w74;
assign w76 = pi041 & ~pi225;
assign w77 = pi043 & ~pi227;
assign w78 = ~w70 & w77;
assign w79 = pi042 & ~pi226;
assign w80 = pi040 & ~pi224;
assign w81 = ~w76 & ~w79;
assign w82 = ~w80 & w81;
assign w83 = ~w78 & w82;
assign w84 = ~w75 & w83;
assign w85 = ~pi039 & pi223;
assign w86 = ~pi040 & pi224;
assign w87 = ~pi041 & pi225;
assign w88 = ~w80 & w87;
assign w89 = ~w86 & ~w88;
assign w90 = ~w85 & w89;
assign w91 = (~w62 & w84) | (~w62 & w16169) | (w84 & w16169);
assign w92 = w61 & w91;
assign w93 = pi046 & ~pi246;
assign w94 = pi045 & ~pi245;
assign w95 = ~w93 & ~w94;
assign w96 = ~pi045 & pi245;
assign w97 = ~pi044 & pi244;
assign w98 = ~w96 & ~w97;
assign w99 = ~w95 & w98;
assign w100 = pi042 & ~pi242;
assign w101 = pi041 & ~pi241;
assign w102 = ~w100 & ~w101;
assign w103 = pi044 & ~pi244;
assign w104 = pi043 & ~pi243;
assign w105 = ~w103 & ~w104;
assign w106 = w102 & w105;
assign w107 = ~w99 & w106;
assign w108 = ~pi043 & pi243;
assign w109 = ~pi042 & pi242;
assign w110 = ~w108 & ~w109;
assign w111 = w102 & ~w110;
assign w112 = ~pi039 & pi239;
assign w113 = ~pi041 & pi241;
assign w114 = ~pi040 & pi240;
assign w115 = ~w113 & ~w114;
assign w116 = ~w112 & w115;
assign w117 = ~w111 & w116;
assign w118 = ~w107 & w117;
assign w119 = pi040 & ~pi240;
assign w120 = pi039 & ~pi239;
assign w121 = ~w119 & ~w120;
assign w122 = ~w112 & ~w121;
assign w123 = ~w118 & ~w122;
assign w124 = pi046 & ~pi238;
assign w125 = pi045 & ~pi237;
assign w126 = ~w124 & ~w125;
assign w127 = ~pi045 & pi237;
assign w128 = ~pi044 & pi236;
assign w129 = ~w127 & ~w128;
assign w130 = ~w126 & w129;
assign w131 = pi042 & ~pi234;
assign w132 = pi041 & ~pi233;
assign w133 = ~w131 & ~w132;
assign w134 = pi044 & ~pi236;
assign w135 = pi043 & ~pi235;
assign w136 = ~w134 & ~w135;
assign w137 = w133 & w136;
assign w138 = ~w130 & w137;
assign w139 = ~pi043 & pi235;
assign w140 = ~pi042 & pi234;
assign w141 = ~w139 & ~w140;
assign w142 = w133 & ~w141;
assign w143 = ~pi039 & pi231;
assign w144 = ~pi041 & pi233;
assign w145 = ~pi040 & pi232;
assign w146 = ~w144 & ~w145;
assign w147 = ~w143 & w146;
assign w148 = ~w142 & w147;
assign w149 = ~w138 & w148;
assign w150 = pi040 & ~pi232;
assign w151 = pi039 & ~pi231;
assign w152 = ~w150 & ~w151;
assign w153 = ~w143 & ~w152;
assign w154 = ~w149 & ~w153;
assign w155 = w123 & w154;
assign w156 = pi046 & ~pi206;
assign w157 = pi045 & ~pi205;
assign w158 = ~w156 & ~w157;
assign w159 = ~pi045 & pi205;
assign w160 = ~pi044 & pi204;
assign w161 = ~w159 & ~w160;
assign w162 = ~w158 & w161;
assign w163 = pi042 & ~pi202;
assign w164 = pi041 & ~pi201;
assign w165 = ~w163 & ~w164;
assign w166 = pi044 & ~pi204;
assign w167 = pi043 & ~pi203;
assign w168 = ~w166 & ~w167;
assign w169 = w165 & w168;
assign w170 = ~w162 & w169;
assign w171 = ~pi043 & pi203;
assign w172 = ~pi042 & pi202;
assign w173 = ~w171 & ~w172;
assign w174 = w165 & ~w173;
assign w175 = ~pi039 & pi199;
assign w176 = ~pi041 & pi201;
assign w177 = ~pi040 & pi200;
assign w178 = ~w176 & ~w177;
assign w179 = ~w175 & w178;
assign w180 = ~w174 & w179;
assign w181 = ~w170 & w180;
assign w182 = pi040 & ~pi200;
assign w183 = pi039 & ~pi199;
assign w184 = ~w182 & ~w183;
assign w185 = ~w175 & ~w184;
assign w186 = ~w181 & ~w185;
assign w187 = pi046 & ~pi214;
assign w188 = pi045 & ~pi213;
assign w189 = ~w187 & ~w188;
assign w190 = ~pi045 & pi213;
assign w191 = ~pi044 & pi212;
assign w192 = ~w190 & ~w191;
assign w193 = ~w189 & w192;
assign w194 = pi042 & ~pi210;
assign w195 = pi041 & ~pi209;
assign w196 = ~w194 & ~w195;
assign w197 = pi044 & ~pi212;
assign w198 = pi043 & ~pi211;
assign w199 = ~w197 & ~w198;
assign w200 = w196 & w199;
assign w201 = ~w193 & w200;
assign w202 = ~pi043 & pi211;
assign w203 = ~pi042 & pi210;
assign w204 = ~w202 & ~w203;
assign w205 = w196 & ~w204;
assign w206 = ~pi039 & pi207;
assign w207 = ~pi041 & pi209;
assign w208 = ~pi040 & pi208;
assign w209 = ~w207 & ~w208;
assign w210 = ~w206 & w209;
assign w211 = ~w205 & w210;
assign w212 = ~w201 & w211;
assign w213 = pi040 & ~pi208;
assign w214 = pi039 & ~pi207;
assign w215 = ~w213 & ~w214;
assign w216 = ~w206 & ~w215;
assign w217 = ~w212 & ~w216;
assign w218 = w186 & w217;
assign w219 = w155 & w218;
assign w220 = w92 & w219;
assign w221 = pi046 & ~pi198;
assign w222 = pi045 & ~pi197;
assign w223 = ~w221 & ~w222;
assign w224 = ~pi045 & pi197;
assign w225 = ~pi044 & pi196;
assign w226 = ~w224 & ~w225;
assign w227 = ~w223 & w226;
assign w228 = pi044 & ~pi196;
assign w229 = pi043 & ~pi195;
assign w230 = ~w228 & ~w229;
assign w231 = ~pi043 & pi195;
assign w232 = ~pi042 & pi194;
assign w233 = ~w231 & ~w232;
assign w234 = (w233 & w227) | (w233 & w16170) | (w227 & w16170);
assign w235 = pi042 & ~pi194;
assign w236 = pi041 & ~pi193;
assign w237 = ~w235 & ~w236;
assign w238 = ~w234 & w237;
assign w239 = ~pi039 & pi191;
assign w240 = ~pi040 & pi192;
assign w241 = ~pi041 & pi193;
assign w242 = ~w239 & ~w240;
assign w243 = ~w241 & w242;
assign w244 = ~w238 & w243;
assign w245 = pi039 & ~pi191;
assign w246 = pi040 & ~pi192;
assign w247 = ~w239 & w246;
assign w248 = ~w245 & ~w247;
assign w249 = ~w244 & w248;
assign w250 = ~pi045 & pi109;
assign w251 = pi046 & ~pi110;
assign w252 = ~w250 & w251;
assign w253 = pi045 & ~pi109;
assign w254 = pi044 & ~pi108;
assign w255 = ~w253 & ~w254;
assign w256 = ~w252 & w255;
assign w257 = ~pi044 & pi108;
assign w258 = ~pi043 & pi107;
assign w259 = ~w257 & ~w258;
assign w260 = pi043 & ~pi107;
assign w261 = pi042 & ~pi106;
assign w262 = ~w260 & ~w261;
assign w263 = (w262 & w256) | (w262 & w16171) | (w256 & w16171);
assign w264 = ~pi042 & pi106;
assign w265 = ~pi041 & pi105;
assign w266 = ~w264 & ~w265;
assign w267 = ~w263 & w266;
assign w268 = pi039 & ~pi103;
assign w269 = pi040 & ~pi104;
assign w270 = pi041 & ~pi105;
assign w271 = ~w268 & ~w269;
assign w272 = ~w270 & w271;
assign w273 = ~w267 & w272;
assign w274 = ~pi039 & pi103;
assign w275 = ~pi040 & pi104;
assign w276 = ~w268 & w275;
assign w277 = ~w274 & ~w276;
assign w278 = ~w273 & w277;
assign w279 = w249 & ~w278;
assign w280 = w220 & w279;
assign w281 = ~pi039 & pi095;
assign w282 = ~pi043 & pi099;
assign w283 = ~pi042 & pi098;
assign w284 = ~w282 & ~w283;
assign w285 = pi044 & ~pi100;
assign w286 = pi043 & ~pi099;
assign w287 = ~w285 & ~w286;
assign w288 = w284 & ~w287;
assign w289 = pi040 & ~pi096;
assign w290 = pi039 & ~pi095;
assign w291 = ~w289 & ~w290;
assign w292 = pi042 & ~pi098;
assign w293 = pi041 & ~pi097;
assign w294 = pi046 & ~pi102;
assign w295 = pi045 & ~pi101;
assign w296 = ~w294 & ~w295;
assign w297 = ~pi045 & pi101;
assign w298 = ~pi044 & pi100;
assign w299 = ~w297 & ~w298;
assign w300 = w284 & w299;
assign w301 = ~w296 & w300;
assign w302 = ~w292 & ~w293;
assign w303 = w291 & w302;
assign w304 = ~w288 & w303;
assign w305 = ~w301 & w304;
assign w306 = ~pi041 & pi097;
assign w307 = ~pi040 & pi096;
assign w308 = ~w306 & ~w307;
assign w309 = w291 & ~w308;
assign w310 = ~w305 & ~w309;
assign w311 = ~w305 & w16172;
assign w312 = pi045 & ~pi093;
assign w313 = pi044 & ~pi092;
assign w314 = ~pi045 & pi093;
assign w315 = pi046 & ~pi094;
assign w316 = ~w314 & w315;
assign w317 = ~w312 & ~w313;
assign w318 = ~w316 & w317;
assign w319 = ~pi044 & pi092;
assign w320 = ~pi042 & pi090;
assign w321 = ~pi041 & pi089;
assign w322 = ~w320 & ~w321;
assign w323 = ~pi043 & pi091;
assign w324 = ~w319 & ~w323;
assign w325 = w322 & w324;
assign w326 = ~w318 & w325;
assign w327 = pi041 & ~pi089;
assign w328 = pi043 & ~pi091;
assign w329 = pi042 & ~pi090;
assign w330 = ~w328 & ~w329;
assign w331 = w322 & ~w330;
assign w332 = pi039 & ~pi087;
assign w333 = pi040 & ~pi088;
assign w334 = ~w327 & ~w332;
assign w335 = ~w333 & w334;
assign w336 = ~w331 & w335;
assign w337 = ~w326 & w336;
assign w338 = ~pi039 & pi087;
assign w339 = ~pi040 & pi088;
assign w340 = ~w332 & w339;
assign w341 = ~w338 & ~w340;
assign w342 = ~w337 & w341;
assign w343 = ~w311 & ~w342;
assign w344 = ~pi039 & pi079;
assign w345 = pi040 & ~pi080;
assign w346 = pi039 & ~pi079;
assign w347 = ~w345 & ~w346;
assign w348 = ~w344 & ~w347;
assign w349 = ~pi043 & pi083;
assign w350 = ~pi042 & pi082;
assign w351 = ~w349 & ~w350;
assign w352 = pi042 & ~pi082;
assign w353 = pi041 & ~pi081;
assign w354 = ~w352 & ~w353;
assign w355 = ~w351 & w354;
assign w356 = pi046 & ~pi086;
assign w357 = pi045 & ~pi085;
assign w358 = ~w356 & ~w357;
assign w359 = ~pi045 & pi085;
assign w360 = ~pi044 & pi084;
assign w361 = ~w359 & ~w360;
assign w362 = ~w358 & w361;
assign w363 = pi044 & ~pi084;
assign w364 = pi043 & ~pi083;
assign w365 = ~w363 & ~w364;
assign w366 = w354 & w365;
assign w367 = ~w362 & w366;
assign w368 = ~pi041 & pi081;
assign w369 = ~pi040 & pi080;
assign w370 = ~w368 & ~w369;
assign w371 = ~w344 & w370;
assign w372 = ~w367 & w16173;
assign w373 = ~w348 & ~w372;
assign w374 = pi045 & ~pi077;
assign w375 = pi044 & ~pi076;
assign w376 = ~pi045 & pi077;
assign w377 = pi046 & ~pi078;
assign w378 = ~w376 & w377;
assign w379 = ~w374 & ~w375;
assign w380 = ~w378 & w379;
assign w381 = ~pi044 & pi076;
assign w382 = ~pi042 & pi074;
assign w383 = ~pi041 & pi073;
assign w384 = ~w382 & ~w383;
assign w385 = ~pi043 & pi075;
assign w386 = ~w381 & ~w385;
assign w387 = w384 & w386;
assign w388 = ~w380 & w387;
assign w389 = pi041 & ~pi073;
assign w390 = pi043 & ~pi075;
assign w391 = pi042 & ~pi074;
assign w392 = ~w390 & ~w391;
assign w393 = w384 & ~w392;
assign w394 = pi039 & ~pi071;
assign w395 = pi040 & ~pi072;
assign w396 = ~w389 & ~w394;
assign w397 = ~w395 & w396;
assign w398 = ~w393 & w397;
assign w399 = ~w388 & w398;
assign w400 = ~pi039 & pi071;
assign w401 = ~pi040 & pi072;
assign w402 = ~w394 & w401;
assign w403 = ~w400 & ~w402;
assign w404 = ~w399 & w403;
assign w405 = w373 & ~w404;
assign w406 = w343 & w405;
assign w407 = ~pi039 & pi063;
assign w408 = ~pi043 & pi067;
assign w409 = ~pi042 & pi066;
assign w410 = ~w408 & ~w409;
assign w411 = pi044 & ~pi068;
assign w412 = pi043 & ~pi067;
assign w413 = ~w411 & ~w412;
assign w414 = w410 & ~w413;
assign w415 = pi040 & ~pi064;
assign w416 = pi039 & ~pi063;
assign w417 = ~w415 & ~w416;
assign w418 = pi042 & ~pi066;
assign w419 = pi041 & ~pi065;
assign w420 = pi046 & ~pi070;
assign w421 = pi045 & ~pi069;
assign w422 = ~w420 & ~w421;
assign w423 = ~pi045 & pi069;
assign w424 = ~pi044 & pi068;
assign w425 = ~w423 & ~w424;
assign w426 = w410 & w425;
assign w427 = ~w422 & w426;
assign w428 = ~w418 & ~w419;
assign w429 = w417 & w428;
assign w430 = ~w414 & w429;
assign w431 = ~w427 & w430;
assign w432 = ~pi041 & pi065;
assign w433 = ~pi040 & pi064;
assign w434 = ~w432 & ~w433;
assign w435 = w417 & ~w434;
assign w436 = ~w431 & ~w435;
assign w437 = ~w407 & w436;
assign w438 = pi043 & ~pi059;
assign w439 = pi044 & ~pi060;
assign w440 = ~pi044 & pi060;
assign w441 = pi046 & ~pi062;
assign w442 = pi045 & ~pi061;
assign w443 = ~w441 & ~w442;
assign w444 = ~pi045 & pi061;
assign w445 = ~w440 & ~w444;
assign w446 = ~w443 & w445;
assign w447 = ~w438 & ~w439;
assign w448 = ~w446 & w447;
assign w449 = ~pi043 & pi059;
assign w450 = ~pi042 & pi058;
assign w451 = ~w449 & ~w450;
assign w452 = ~w448 & w451;
assign w453 = pi042 & ~pi058;
assign w454 = pi040 & ~pi056;
assign w455 = pi039 & ~pi055;
assign w456 = ~w454 & ~w455;
assign w457 = pi041 & ~pi057;
assign w458 = ~w453 & ~w457;
assign w459 = w456 & w458;
assign w460 = ~w452 & w459;
assign w461 = ~pi039 & pi055;
assign w462 = ~pi041 & pi057;
assign w463 = ~pi040 & pi056;
assign w464 = ~w462 & ~w463;
assign w465 = w456 & ~w464;
assign w466 = ~w461 & ~w465;
assign w467 = ~w460 & w466;
assign w468 = ~w437 & ~w467;
assign w469 = w406 & w468;
assign w470 = w280 & w469;
assign w471 = ~pi039 & pi247;
assign w472 = pi040 & ~pi248;
assign w473 = pi039 & ~pi247;
assign w474 = ~w472 & ~w473;
assign w475 = ~w471 & ~w474;
assign w476 = ~pi043 & pi251;
assign w477 = ~pi042 & pi250;
assign w478 = ~w476 & ~w477;
assign w479 = pi042 & ~pi250;
assign w480 = pi041 & ~pi249;
assign w481 = ~w479 & ~w480;
assign w482 = ~w478 & w481;
assign w483 = pi046 & ~pi254;
assign w484 = pi045 & ~pi253;
assign w485 = ~w483 & ~w484;
assign w486 = ~pi045 & pi253;
assign w487 = ~pi044 & pi252;
assign w488 = ~w486 & ~w487;
assign w489 = ~w485 & w488;
assign w490 = pi044 & ~pi252;
assign w491 = pi043 & ~pi251;
assign w492 = ~w490 & ~w491;
assign w493 = w481 & w492;
assign w494 = ~w489 & w493;
assign w495 = ~w482 & ~w494;
assign w496 = ~pi041 & pi249;
assign w497 = ~pi040 & pi248;
assign w498 = ~w496 & ~w497;
assign w499 = ~w471 & w498;
assign w500 = ~w494 & w16174;
assign w501 = ~w475 & ~w500;
assign w502 = pi046 & ~pi262;
assign w503 = pi045 & ~pi261;
assign w504 = ~w502 & ~w503;
assign w505 = ~pi045 & pi261;
assign w506 = ~pi044 & pi260;
assign w507 = ~w505 & ~w506;
assign w508 = ~w504 & w507;
assign w509 = pi044 & ~pi260;
assign w510 = pi043 & ~pi259;
assign w511 = ~w509 & ~w510;
assign w512 = ~w508 & w511;
assign w513 = pi040 & ~pi256;
assign w514 = pi039 & ~pi255;
assign w515 = ~w513 & ~w514;
assign w516 = ~pi041 & pi257;
assign w517 = ~pi040 & pi256;
assign w518 = ~w516 & ~w517;
assign w519 = w515 & ~w518;
assign w520 = ~pi043 & pi259;
assign w521 = ~pi042 & pi258;
assign w522 = ~w520 & ~w521;
assign w523 = ~w519 & w522;
assign w524 = ~w512 & w523;
assign w525 = pi042 & ~pi258;
assign w526 = pi041 & ~pi257;
assign w527 = ~w525 & ~w526;
assign w528 = w518 & ~w527;
assign w529 = w515 & ~w528;
assign w530 = ~w524 & w529;
assign w531 = ~pi039 & pi255;
assign w532 = (~w531 & w524) | (~w531 & w16175) | (w524 & w16175);
assign w533 = w501 & ~w532;
assign w534 = ~pi043 & pi275;
assign w535 = ~pi042 & pi274;
assign w536 = ~w534 & ~w535;
assign w537 = pi044 & ~pi276;
assign w538 = pi043 & ~pi275;
assign w539 = ~w537 & ~w538;
assign w540 = w536 & ~w539;
assign w541 = pi040 & ~pi272;
assign w542 = pi039 & ~pi271;
assign w543 = ~w541 & ~w542;
assign w544 = pi042 & ~pi274;
assign w545 = pi041 & ~pi273;
assign w546 = pi046 & ~pi278;
assign w547 = pi045 & ~pi277;
assign w548 = ~w546 & ~w547;
assign w549 = ~pi045 & pi277;
assign w550 = ~pi044 & pi276;
assign w551 = ~w549 & ~w550;
assign w552 = w536 & w551;
assign w553 = ~w548 & w552;
assign w554 = ~w544 & ~w545;
assign w555 = w543 & w554;
assign w556 = ~w540 & w555;
assign w557 = ~w553 & w556;
assign w558 = ~pi041 & pi273;
assign w559 = ~pi040 & pi272;
assign w560 = ~w558 & ~w559;
assign w561 = w543 & ~w560;
assign w562 = ~w557 & ~w561;
assign w563 = ~pi039 & pi271;
assign w564 = ~w557 & w16176;
assign w565 = ~pi043 & pi267;
assign w566 = ~pi042 & pi266;
assign w567 = ~w565 & ~w566;
assign w568 = pi044 & ~pi268;
assign w569 = pi043 & ~pi267;
assign w570 = ~w568 & ~w569;
assign w571 = w567 & ~w570;
assign w572 = pi040 & ~pi264;
assign w573 = pi039 & ~pi263;
assign w574 = ~w572 & ~w573;
assign w575 = pi042 & ~pi266;
assign w576 = pi041 & ~pi265;
assign w577 = pi046 & ~pi270;
assign w578 = pi045 & ~pi269;
assign w579 = ~w577 & ~w578;
assign w580 = ~pi045 & pi269;
assign w581 = ~pi044 & pi268;
assign w582 = ~w580 & ~w581;
assign w583 = w567 & w582;
assign w584 = ~w579 & w583;
assign w585 = ~w575 & ~w576;
assign w586 = w574 & w585;
assign w587 = ~w571 & w586;
assign w588 = ~w584 & w587;
assign w589 = ~pi041 & pi265;
assign w590 = ~pi040 & pi264;
assign w591 = ~w589 & ~w590;
assign w592 = w574 & ~w591;
assign w593 = ~w588 & ~w592;
assign w594 = ~pi039 & pi263;
assign w595 = ~w588 & w16177;
assign w596 = ~w564 & ~w595;
assign w597 = w533 & w596;
assign w598 = pi046 & ~pi174;
assign w599 = pi045 & ~pi173;
assign w600 = ~w598 & ~w599;
assign w601 = ~pi045 & pi173;
assign w602 = ~pi044 & pi172;
assign w603 = ~w601 & ~w602;
assign w604 = ~w600 & w603;
assign w605 = pi042 & ~pi170;
assign w606 = pi041 & ~pi169;
assign w607 = ~w605 & ~w606;
assign w608 = pi044 & ~pi172;
assign w609 = pi043 & ~pi171;
assign w610 = ~w608 & ~w609;
assign w611 = w607 & w610;
assign w612 = ~w604 & w611;
assign w613 = ~pi043 & pi171;
assign w614 = ~pi042 & pi170;
assign w615 = ~w613 & ~w614;
assign w616 = w607 & ~w615;
assign w617 = ~pi039 & pi167;
assign w618 = ~pi041 & pi169;
assign w619 = ~pi040 & pi168;
assign w620 = ~w618 & ~w619;
assign w621 = ~w617 & w620;
assign w622 = ~w616 & w621;
assign w623 = ~w612 & w622;
assign w624 = pi040 & ~pi168;
assign w625 = pi039 & ~pi167;
assign w626 = ~w624 & ~w625;
assign w627 = ~w617 & ~w626;
assign w628 = ~w623 & ~w627;
assign w629 = ~pi045 & pi181;
assign w630 = pi046 & ~pi182;
assign w631 = ~w629 & w630;
assign w632 = pi045 & ~pi181;
assign w633 = pi044 & ~pi180;
assign w634 = ~w632 & ~w633;
assign w635 = ~w631 & w634;
assign w636 = ~pi042 & pi178;
assign w637 = ~pi041 & pi177;
assign w638 = ~w636 & ~w637;
assign w639 = ~pi044 & pi180;
assign w640 = ~pi043 & pi179;
assign w641 = ~w639 & ~w640;
assign w642 = w638 & w641;
assign w643 = ~w635 & w642;
assign w644 = pi043 & ~pi179;
assign w645 = pi042 & ~pi178;
assign w646 = ~w644 & ~w645;
assign w647 = w638 & ~w646;
assign w648 = pi041 & ~pi177;
assign w649 = pi039 & ~pi175;
assign w650 = pi040 & ~pi176;
assign w651 = ~w648 & ~w649;
assign w652 = ~w650 & w651;
assign w653 = ~w647 & w652;
assign w654 = ~w643 & w653;
assign w655 = ~pi039 & pi175;
assign w656 = ~pi040 & pi176;
assign w657 = ~w649 & w656;
assign w658 = ~w655 & ~w657;
assign w659 = ~w654 & w658;
assign w660 = w628 & ~w659;
assign w661 = pi043 & ~pi163;
assign w662 = pi044 & ~pi164;
assign w663 = ~pi044 & pi164;
assign w664 = pi046 & ~pi166;
assign w665 = pi045 & ~pi165;
assign w666 = ~w664 & ~w665;
assign w667 = ~pi045 & pi165;
assign w668 = ~w663 & ~w667;
assign w669 = ~w666 & w668;
assign w670 = ~w661 & ~w662;
assign w671 = ~w669 & w670;
assign w672 = ~pi042 & pi162;
assign w673 = ~pi043 & pi163;
assign w674 = ~pi041 & pi161;
assign w675 = ~pi039 & pi159;
assign w676 = ~pi040 & pi160;
assign w677 = ~w674 & ~w675;
assign w678 = ~w676 & w677;
assign w679 = ~w672 & ~w673;
assign w680 = w678 & w679;
assign w681 = ~w671 & w680;
assign w682 = pi039 & ~pi159;
assign w683 = pi042 & ~pi162;
assign w684 = pi041 & ~pi161;
assign w685 = ~w683 & ~w684;
assign w686 = w678 & ~w685;
assign w687 = pi040 & ~pi160;
assign w688 = ~w675 & w687;
assign w689 = ~w682 & ~w688;
assign w690 = ~w686 & w689;
assign w691 = ~w681 & w690;
assign w692 = w660 & w691;
assign w693 = ~pi039 & pi111;
assign w694 = pi040 & ~pi112;
assign w695 = pi039 & ~pi111;
assign w696 = ~w694 & ~w695;
assign w697 = ~w693 & ~w696;
assign w698 = ~pi043 & pi115;
assign w699 = ~pi042 & pi114;
assign w700 = ~w698 & ~w699;
assign w701 = pi042 & ~pi114;
assign w702 = pi041 & ~pi113;
assign w703 = ~w701 & ~w702;
assign w704 = ~w700 & w703;
assign w705 = pi046 & ~pi118;
assign w706 = pi045 & ~pi117;
assign w707 = ~w705 & ~w706;
assign w708 = ~pi045 & pi117;
assign w709 = ~pi044 & pi116;
assign w710 = ~w708 & ~w709;
assign w711 = ~w707 & w710;
assign w712 = pi044 & ~pi116;
assign w713 = pi043 & ~pi115;
assign w714 = ~w712 & ~w713;
assign w715 = w703 & w714;
assign w716 = ~w711 & w715;
assign w717 = ~w704 & ~w716;
assign w718 = ~pi041 & pi113;
assign w719 = ~pi040 & pi112;
assign w720 = ~w718 & ~w719;
assign w721 = ~w693 & w720;
assign w722 = ~w716 & w16178;
assign w723 = ~w697 & ~w722;
assign w724 = pi043 & ~pi123;
assign w725 = pi044 & ~pi124;
assign w726 = ~pi044 & pi124;
assign w727 = pi046 & ~pi126;
assign w728 = pi045 & ~pi125;
assign w729 = ~w727 & ~w728;
assign w730 = ~pi045 & pi125;
assign w731 = ~w726 & ~w730;
assign w732 = ~w729 & w731;
assign w733 = ~w724 & ~w725;
assign w734 = ~w732 & w733;
assign w735 = ~pi042 & pi122;
assign w736 = ~pi043 & pi123;
assign w737 = ~pi041 & pi121;
assign w738 = ~pi039 & pi119;
assign w739 = ~pi040 & pi120;
assign w740 = ~w737 & ~w738;
assign w741 = ~w739 & w740;
assign w742 = ~w735 & ~w736;
assign w743 = w741 & w742;
assign w744 = ~w734 & w743;
assign w745 = pi039 & ~pi119;
assign w746 = pi042 & ~pi122;
assign w747 = pi041 & ~pi121;
assign w748 = ~w746 & ~w747;
assign w749 = w741 & ~w748;
assign w750 = pi040 & ~pi120;
assign w751 = ~w738 & w750;
assign w752 = ~w745 & ~w751;
assign w753 = ~w749 & w752;
assign w754 = ~w744 & w753;
assign w755 = w723 & w754;
assign w756 = w692 & w755;
assign w757 = w597 & w756;
assign w758 = ~pi045 & pi157;
assign w759 = pi046 & ~pi158;
assign w760 = ~w758 & w759;
assign w761 = pi045 & ~pi157;
assign w762 = pi156 & ~w761;
assign w763 = ~w760 & w762;
assign w764 = pi044 & ~w763;
assign w765 = pi043 & ~pi155;
assign w766 = ~w761 & ~w765;
assign w767 = ~w760 & w766;
assign w768 = pi156 & ~w765;
assign w769 = ~w767 & ~w768;
assign w770 = ~w764 & ~w769;
assign w771 = ~pi042 & pi154;
assign w772 = ~pi041 & pi153;
assign w773 = ~pi040 & pi152;
assign w774 = ~w772 & ~w773;
assign w775 = pi040 & ~pi152;
assign w776 = pi039 & ~pi151;
assign w777 = ~w775 & ~w776;
assign w778 = ~w774 & w777;
assign w779 = ~pi043 & pi155;
assign w780 = ~w771 & ~w779;
assign w781 = ~w778 & w780;
assign w782 = pi042 & ~pi154;
assign w783 = pi041 & ~pi153;
assign w784 = ~w782 & ~w783;
assign w785 = w774 & ~w784;
assign w786 = w777 & ~w785;
assign w787 = (w786 & w770) | (w786 & w16179) | (w770 & w16179);
assign w788 = ~pi039 & pi151;
assign w789 = ~w787 & ~w788;
assign w790 = ~pi045 & pi189;
assign w791 = pi046 & ~pi190;
assign w792 = ~w790 & w791;
assign w793 = pi045 & ~pi189;
assign w794 = pi188 & ~w793;
assign w795 = ~w792 & w794;
assign w796 = pi044 & ~w795;
assign w797 = pi043 & ~pi187;
assign w798 = ~w793 & ~w797;
assign w799 = ~w792 & w798;
assign w800 = pi188 & ~w797;
assign w801 = ~w799 & ~w800;
assign w802 = ~w796 & ~w801;
assign w803 = ~pi042 & pi186;
assign w804 = ~pi041 & pi185;
assign w805 = ~pi040 & pi184;
assign w806 = ~w804 & ~w805;
assign w807 = pi040 & ~pi184;
assign w808 = pi039 & ~pi183;
assign w809 = ~w807 & ~w808;
assign w810 = ~w806 & w809;
assign w811 = ~pi043 & pi187;
assign w812 = ~w803 & ~w811;
assign w813 = ~w810 & w812;
assign w814 = pi042 & ~pi186;
assign w815 = pi041 & ~pi185;
assign w816 = ~w814 & ~w815;
assign w817 = w806 & ~w816;
assign w818 = w809 & ~w817;
assign w819 = (w818 & w802) | (w818 & w16180) | (w802 & w16180);
assign w820 = ~pi039 & pi183;
assign w821 = ~w819 & ~w820;
assign w822 = ~w789 & ~w821;
assign w823 = ~pi039 & pi127;
assign w824 = ~pi040 & pi128;
assign w825 = ~pi045 & pi133;
assign w826 = pi046 & ~pi134;
assign w827 = ~w825 & w826;
assign w828 = pi045 & ~pi133;
assign w829 = pi044 & ~pi132;
assign w830 = ~w828 & ~w829;
assign w831 = ~w827 & w830;
assign w832 = ~pi042 & pi130;
assign w833 = ~pi041 & pi129;
assign w834 = ~w832 & ~w833;
assign w835 = ~pi044 & pi132;
assign w836 = ~pi043 & pi131;
assign w837 = ~w835 & ~w836;
assign w838 = w834 & w837;
assign w839 = ~w831 & w838;
assign w840 = pi043 & ~pi131;
assign w841 = pi042 & ~pi130;
assign w842 = ~w840 & ~w841;
assign w843 = w834 & ~w842;
assign w844 = pi041 & ~pi129;
assign w845 = pi040 & ~pi128;
assign w846 = ~w844 & ~w845;
assign w847 = ~w843 & w846;
assign w848 = ~w839 & w847;
assign w849 = ~w824 & ~w848;
assign w850 = pi039 & ~pi127;
assign w851 = (~w850 & w848) | (~w850 & w16181) | (w848 & w16181);
assign w852 = ~w823 & ~w851;
assign w853 = pi045 & ~pi149;
assign w854 = pi044 & ~pi148;
assign w855 = ~pi045 & pi149;
assign w856 = pi046 & ~pi150;
assign w857 = ~w855 & w856;
assign w858 = ~w853 & ~w854;
assign w859 = ~w857 & w858;
assign w860 = ~pi044 & pi148;
assign w861 = ~pi042 & pi146;
assign w862 = ~pi041 & pi145;
assign w863 = ~w861 & ~w862;
assign w864 = ~pi043 & pi147;
assign w865 = ~w860 & ~w864;
assign w866 = w863 & w865;
assign w867 = ~w859 & w866;
assign w868 = pi039 & ~pi143;
assign w869 = pi043 & ~pi147;
assign w870 = pi042 & ~pi146;
assign w871 = ~w869 & ~w870;
assign w872 = w863 & ~w871;
assign w873 = pi040 & ~pi144;
assign w874 = pi041 & ~pi145;
assign w875 = ~w868 & ~w873;
assign w876 = ~w874 & w875;
assign w877 = ~w872 & w876;
assign w878 = ~w867 & w877;
assign w879 = ~pi039 & pi143;
assign w880 = ~pi040 & pi144;
assign w881 = ~w868 & w880;
assign w882 = ~w879 & ~w881;
assign w883 = ~w878 & w882;
assign w884 = pi039 & ~pi135;
assign w885 = ~pi043 & pi139;
assign w886 = ~pi042 & pi138;
assign w887 = ~w885 & ~w886;
assign w888 = pi044 & ~pi140;
assign w889 = pi043 & ~pi139;
assign w890 = ~w888 & ~w889;
assign w891 = w887 & ~w890;
assign w892 = pi041 & ~pi137;
assign w893 = pi040 & ~pi136;
assign w894 = pi042 & ~pi138;
assign w895 = pi046 & ~pi142;
assign w896 = pi045 & ~pi141;
assign w897 = ~w895 & ~w896;
assign w898 = ~pi045 & pi141;
assign w899 = ~pi044 & pi140;
assign w900 = ~w898 & ~w899;
assign w901 = w887 & w900;
assign w902 = ~w897 & w901;
assign w903 = ~w892 & ~w893;
assign w904 = ~w894 & w903;
assign w905 = ~w891 & w904;
assign w906 = ~w902 & w905;
assign w907 = ~pi039 & pi135;
assign w908 = ~pi040 & pi136;
assign w909 = ~pi041 & pi137;
assign w910 = ~w893 & w909;
assign w911 = ~w908 & ~w910;
assign w912 = ~w907 & w911;
assign w913 = (~w884 & w906) | (~w884 & w16182) | (w906 & w16182);
assign w914 = ~w883 & w913;
assign w915 = ~w852 & w914;
assign w916 = w822 & w915;
assign w917 = w757 & w916;
assign w918 = w470 & w917;
assign w919 = ~w29 & w918;
assign w920 = pi001 & w919;
assign w921 = ~w30 & ~w920;
assign w922 = ~w27 & w436;
assign w923 = pi062 & ~pi070;
assign w924 = pi061 & ~pi069;
assign w925 = ~w923 & ~w924;
assign w926 = ~pi061 & pi069;
assign w927 = ~pi060 & pi068;
assign w928 = ~w926 & ~w927;
assign w929 = ~w925 & w928;
assign w930 = pi060 & ~pi068;
assign w931 = pi059 & ~pi067;
assign w932 = ~w930 & ~w931;
assign w933 = ~w929 & w932;
assign w934 = ~pi058 & pi066;
assign w935 = ~pi057 & pi065;
assign w936 = ~pi056 & pi064;
assign w937 = ~w935 & ~w936;
assign w938 = ~pi059 & pi067;
assign w939 = ~w934 & ~w938;
assign w940 = w937 & w939;
assign w941 = ~w933 & w940;
assign w942 = pi056 & ~pi064;
assign w943 = pi058 & ~pi066;
assign w944 = pi057 & ~pi065;
assign w945 = ~w943 & ~w944;
assign w946 = w937 & ~w945;
assign w947 = pi055 & ~pi063;
assign w948 = ~w942 & ~w947;
assign w949 = ~w946 & w948;
assign w950 = ~w941 & w949;
assign w951 = ~pi055 & pi063;
assign w952 = ~w28 & ~w407;
assign w953 = ~w951 & w952;
assign w954 = (w953 & w941) | (w953 & w16183) | (w941 & w16183);
assign w955 = w922 & w954;
assign w956 = pi004 & w955;
assign w957 = ~pi055 & pi095;
assign w958 = pi062 & ~pi102;
assign w959 = pi061 & ~pi101;
assign w960 = ~w958 & ~w959;
assign w961 = ~pi061 & pi101;
assign w962 = ~pi060 & pi100;
assign w963 = ~w961 & ~w962;
assign w964 = ~w960 & w963;
assign w965 = pi060 & ~pi100;
assign w966 = pi059 & ~pi099;
assign w967 = ~w965 & ~w966;
assign w968 = ~pi059 & pi099;
assign w969 = ~pi058 & pi098;
assign w970 = ~w968 & ~w969;
assign w971 = (w970 & w964) | (w970 & w16184) | (w964 & w16184);
assign w972 = pi058 & ~pi098;
assign w973 = pi057 & ~pi097;
assign w974 = ~w972 & ~w973;
assign w975 = ~w971 & w974;
assign w976 = ~pi057 & pi097;
assign w977 = ~pi056 & pi096;
assign w978 = ~w976 & ~w977;
assign w979 = ~w975 & w978;
assign w980 = pi056 & ~pi096;
assign w981 = pi055 & ~pi095;
assign w982 = ~w980 & ~w981;
assign w983 = ~w979 & w982;
assign w984 = ~w957 & ~w983;
assign w985 = pi055 & ~pi087;
assign w986 = ~pi061 & pi093;
assign w987 = pi062 & ~pi094;
assign w988 = ~w986 & w987;
assign w989 = pi061 & ~pi093;
assign w990 = pi060 & ~pi092;
assign w991 = ~w989 & ~w990;
assign w992 = ~w988 & w991;
assign w993 = ~pi060 & pi092;
assign w994 = ~pi059 & pi091;
assign w995 = ~w993 & ~w994;
assign w996 = pi059 & ~pi091;
assign w997 = pi058 & ~pi090;
assign w998 = ~w996 & ~w997;
assign w999 = (w998 & w992) | (w998 & w16185) | (w992 & w16185);
assign w1000 = ~pi058 & pi090;
assign w1001 = ~pi057 & pi089;
assign w1002 = ~w1000 & ~w1001;
assign w1003 = ~w999 & w1002;
assign w1004 = pi056 & ~pi088;
assign w1005 = pi057 & ~pi089;
assign w1006 = ~w1004 & ~w1005;
assign w1007 = ~w1003 & w1006;
assign w1008 = ~pi055 & pi087;
assign w1009 = ~pi056 & pi088;
assign w1010 = ~w1008 & ~w1009;
assign w1011 = ~w1007 & w1010;
assign w1012 = ~w985 & ~w1011;
assign w1013 = ~w984 & w1012;
assign w1014 = ~pi055 & pi135;
assign w1015 = ~pi061 & pi141;
assign w1016 = pi062 & ~pi142;
assign w1017 = pi061 & ~pi141;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = ~pi060 & pi140;
assign w1020 = ~w1015 & ~w1019;
assign w1021 = ~w1018 & w1020;
assign w1022 = pi059 & ~pi139;
assign w1023 = pi058 & ~pi138;
assign w1024 = pi057 & ~pi137;
assign w1025 = ~w1023 & ~w1024;
assign w1026 = pi060 & ~pi140;
assign w1027 = ~w1022 & ~w1026;
assign w1028 = w1025 & w1027;
assign w1029 = ~w1021 & w1028;
assign w1030 = ~pi056 & pi136;
assign w1031 = ~pi059 & pi139;
assign w1032 = ~pi058 & pi138;
assign w1033 = ~w1031 & ~w1032;
assign w1034 = w1025 & ~w1033;
assign w1035 = ~pi057 & pi137;
assign w1036 = ~w1030 & ~w1035;
assign w1037 = ~w1034 & w1036;
assign w1038 = ~w1029 & w1037;
assign w1039 = pi056 & ~pi136;
assign w1040 = pi055 & ~pi135;
assign w1041 = ~w1039 & ~w1040;
assign w1042 = ~w1038 & w1041;
assign w1043 = (~w1014 & w1038) | (~w1014 & w16186) | (w1038 & w16186);
assign w1044 = pi062 & ~pi174;
assign w1045 = pi061 & ~pi173;
assign w1046 = ~w1044 & ~w1045;
assign w1047 = ~pi061 & pi173;
assign w1048 = ~pi060 & pi172;
assign w1049 = ~w1047 & ~w1048;
assign w1050 = ~w1046 & w1049;
assign w1051 = pi058 & ~pi170;
assign w1052 = pi057 & ~pi169;
assign w1053 = ~w1051 & ~w1052;
assign w1054 = pi060 & ~pi172;
assign w1055 = pi059 & ~pi171;
assign w1056 = ~w1054 & ~w1055;
assign w1057 = w1053 & w1056;
assign w1058 = ~w1050 & w1057;
assign w1059 = ~pi059 & pi171;
assign w1060 = ~pi058 & pi170;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = w1053 & ~w1061;
assign w1063 = ~pi057 & pi169;
assign w1064 = ~pi056 & pi168;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = ~w1062 & w1065;
assign w1067 = ~w1058 & w1066;
assign w1068 = pi056 & ~pi168;
assign w1069 = pi055 & ~pi167;
assign w1070 = ~w1068 & ~w1069;
assign w1071 = ~w1067 & w1070;
assign w1072 = ~pi055 & pi167;
assign w1073 = ~w1071 & ~w1072;
assign w1074 = pi061 & ~pi149;
assign w1075 = pi060 & ~pi148;
assign w1076 = ~pi061 & pi149;
assign w1077 = pi062 & ~pi150;
assign w1078 = ~w1076 & w1077;
assign w1079 = ~w1074 & ~w1075;
assign w1080 = ~w1078 & w1079;
assign w1081 = ~pi060 & pi148;
assign w1082 = ~pi058 & pi146;
assign w1083 = ~pi057 & pi145;
assign w1084 = ~w1082 & ~w1083;
assign w1085 = ~pi059 & pi147;
assign w1086 = ~w1081 & ~w1085;
assign w1087 = w1084 & w1086;
assign w1088 = ~w1080 & w1087;
assign w1089 = pi057 & ~pi145;
assign w1090 = pi059 & ~pi147;
assign w1091 = pi058 & ~pi146;
assign w1092 = ~w1090 & ~w1091;
assign w1093 = w1084 & ~w1092;
assign w1094 = pi055 & ~pi143;
assign w1095 = pi056 & ~pi144;
assign w1096 = ~w1089 & ~w1094;
assign w1097 = ~w1095 & w1096;
assign w1098 = ~w1093 & w1097;
assign w1099 = ~w1088 & w1098;
assign w1100 = ~pi055 & pi143;
assign w1101 = ~pi056 & pi144;
assign w1102 = ~w1094 & w1101;
assign w1103 = ~w1100 & ~w1102;
assign w1104 = ~w1099 & w1103;
assign w1105 = ~w1043 & ~w1104;
assign w1106 = ~w1073 & w1105;
assign w1107 = ~pi061 & pi181;
assign w1108 = pi062 & ~pi182;
assign w1109 = ~w1107 & w1108;
assign w1110 = pi061 & ~pi181;
assign w1111 = pi060 & ~pi180;
assign w1112 = ~w1110 & ~w1111;
assign w1113 = ~w1109 & w1112;
assign w1114 = ~pi058 & pi178;
assign w1115 = ~pi057 & pi177;
assign w1116 = ~w1114 & ~w1115;
assign w1117 = ~pi060 & pi180;
assign w1118 = ~pi059 & pi179;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = w1116 & w1119;
assign w1121 = ~w1113 & w1120;
assign w1122 = pi059 & ~pi179;
assign w1123 = pi058 & ~pi178;
assign w1124 = ~w1122 & ~w1123;
assign w1125 = w1116 & ~w1124;
assign w1126 = pi056 & ~pi176;
assign w1127 = pi055 & ~pi175;
assign w1128 = pi057 & ~pi177;
assign w1129 = ~w1126 & ~w1127;
assign w1130 = ~w1128 & w1129;
assign w1131 = ~w1125 & w1130;
assign w1132 = ~w1121 & w1131;
assign w1133 = ~pi055 & pi175;
assign w1134 = ~pi056 & pi176;
assign w1135 = ~w1127 & w1134;
assign w1136 = ~w1133 & ~w1135;
assign w1137 = ~w1132 & w1136;
assign w1138 = ~pi061 & pi197;
assign w1139 = pi062 & ~pi198;
assign w1140 = ~w1138 & w1139;
assign w1141 = pi061 & ~pi197;
assign w1142 = pi060 & ~pi196;
assign w1143 = ~w1141 & ~w1142;
assign w1144 = ~w1140 & w1143;
assign w1145 = ~pi058 & pi194;
assign w1146 = ~pi057 & pi193;
assign w1147 = ~w1145 & ~w1146;
assign w1148 = ~pi060 & pi196;
assign w1149 = ~pi059 & pi195;
assign w1150 = ~w1148 & ~w1149;
assign w1151 = w1147 & w1150;
assign w1152 = ~w1144 & w1151;
assign w1153 = pi059 & ~pi195;
assign w1154 = pi058 & ~pi194;
assign w1155 = ~w1153 & ~w1154;
assign w1156 = w1147 & ~w1155;
assign w1157 = pi056 & ~pi192;
assign w1158 = pi055 & ~pi191;
assign w1159 = pi057 & ~pi193;
assign w1160 = ~w1157 & ~w1158;
assign w1161 = ~w1159 & w1160;
assign w1162 = ~w1156 & w1161;
assign w1163 = ~w1152 & w1162;
assign w1164 = ~pi055 & pi191;
assign w1165 = ~pi056 & pi192;
assign w1166 = ~w1158 & w1165;
assign w1167 = ~w1164 & ~w1166;
assign w1168 = ~w1163 & w1167;
assign w1169 = ~w1137 & ~w1168;
assign w1170 = ~pi055 & pi079;
assign w1171 = pi062 & ~pi086;
assign w1172 = pi061 & ~pi085;
assign w1173 = ~w1171 & ~w1172;
assign w1174 = ~pi061 & pi085;
assign w1175 = ~pi060 & pi084;
assign w1176 = ~w1174 & ~w1175;
assign w1177 = ~w1173 & w1176;
assign w1178 = pi058 & ~pi082;
assign w1179 = pi057 & ~pi081;
assign w1180 = ~w1178 & ~w1179;
assign w1181 = pi060 & ~pi084;
assign w1182 = pi059 & ~pi083;
assign w1183 = ~w1181 & ~w1182;
assign w1184 = w1180 & w1183;
assign w1185 = ~w1177 & w1184;
assign w1186 = ~pi059 & pi083;
assign w1187 = ~pi058 & pi082;
assign w1188 = ~w1186 & ~w1187;
assign w1189 = w1180 & ~w1188;
assign w1190 = ~pi057 & pi081;
assign w1191 = ~pi056 & pi080;
assign w1192 = ~w1190 & ~w1191;
assign w1193 = ~w1189 & w1192;
assign w1194 = ~w1185 & w1193;
assign w1195 = pi056 & ~pi080;
assign w1196 = pi055 & ~pi079;
assign w1197 = ~w1195 & ~w1196;
assign w1198 = ~w1194 & w1197;
assign w1199 = (~w1170 & w1194) | (~w1170 & w16187) | (w1194 & w16187);
assign w1200 = pi061 & ~pi077;
assign w1201 = pi060 & ~pi076;
assign w1202 = ~pi061 & pi077;
assign w1203 = pi062 & ~pi078;
assign w1204 = ~w1202 & w1203;
assign w1205 = ~w1200 & ~w1201;
assign w1206 = ~w1204 & w1205;
assign w1207 = ~pi060 & pi076;
assign w1208 = ~pi058 & pi074;
assign w1209 = ~pi057 & pi073;
assign w1210 = ~w1208 & ~w1209;
assign w1211 = ~pi059 & pi075;
assign w1212 = ~w1207 & ~w1211;
assign w1213 = w1210 & w1212;
assign w1214 = ~w1206 & w1213;
assign w1215 = pi055 & ~pi071;
assign w1216 = pi059 & ~pi075;
assign w1217 = pi058 & ~pi074;
assign w1218 = ~w1216 & ~w1217;
assign w1219 = w1210 & ~w1218;
assign w1220 = pi056 & ~pi072;
assign w1221 = pi057 & ~pi073;
assign w1222 = ~w1215 & ~w1220;
assign w1223 = ~w1221 & w1222;
assign w1224 = ~w1219 & w1223;
assign w1225 = ~w1214 & w1224;
assign w1226 = ~pi055 & pi071;
assign w1227 = ~pi056 & pi072;
assign w1228 = ~w1215 & w1227;
assign w1229 = ~w1226 & ~w1228;
assign w1230 = ~w1225 & w1229;
assign w1231 = pi062 & ~pi134;
assign w1232 = pi061 & ~pi133;
assign w1233 = ~w1231 & ~w1232;
assign w1234 = ~pi061 & pi133;
assign w1235 = ~pi060 & pi132;
assign w1236 = ~w1234 & ~w1235;
assign w1237 = ~w1233 & w1236;
assign w1238 = pi058 & ~pi130;
assign w1239 = pi057 & ~pi129;
assign w1240 = ~w1238 & ~w1239;
assign w1241 = pi060 & ~pi132;
assign w1242 = pi059 & ~pi131;
assign w1243 = ~w1241 & ~w1242;
assign w1244 = w1240 & w1243;
assign w1245 = ~w1237 & w1244;
assign w1246 = ~pi059 & pi131;
assign w1247 = ~pi058 & pi130;
assign w1248 = ~w1246 & ~w1247;
assign w1249 = w1240 & ~w1248;
assign w1250 = ~pi055 & pi127;
assign w1251 = ~pi057 & pi129;
assign w1252 = ~pi056 & pi128;
assign w1253 = ~w1251 & ~w1252;
assign w1254 = ~w1250 & w1253;
assign w1255 = ~w1249 & w1254;
assign w1256 = ~w1245 & w1255;
assign w1257 = pi056 & ~pi128;
assign w1258 = pi055 & ~pi127;
assign w1259 = ~w1257 & ~w1258;
assign w1260 = ~w1250 & ~w1259;
assign w1261 = ~w1256 & ~w1260;
assign w1262 = ~pi061 & pi125;
assign w1263 = pi062 & ~pi126;
assign w1264 = ~w1262 & w1263;
assign w1265 = pi061 & ~pi125;
assign w1266 = pi060 & ~pi124;
assign w1267 = ~w1265 & ~w1266;
assign w1268 = ~w1264 & w1267;
assign w1269 = ~pi058 & pi122;
assign w1270 = ~pi057 & pi121;
assign w1271 = ~w1269 & ~w1270;
assign w1272 = ~pi060 & pi124;
assign w1273 = ~pi059 & pi123;
assign w1274 = ~w1272 & ~w1273;
assign w1275 = w1271 & w1274;
assign w1276 = ~w1268 & w1275;
assign w1277 = pi059 & ~pi123;
assign w1278 = pi058 & ~pi122;
assign w1279 = ~w1277 & ~w1278;
assign w1280 = w1271 & ~w1279;
assign w1281 = pi057 & ~pi121;
assign w1282 = pi055 & ~pi119;
assign w1283 = pi056 & ~pi120;
assign w1284 = ~w1281 & ~w1282;
assign w1285 = ~w1283 & w1284;
assign w1286 = ~w1280 & w1285;
assign w1287 = ~w1276 & w1286;
assign w1288 = ~pi055 & pi119;
assign w1289 = ~pi056 & pi120;
assign w1290 = ~w1282 & w1289;
assign w1291 = ~w1288 & ~w1290;
assign w1292 = ~w1287 & w1291;
assign w1293 = w1261 & ~w1292;
assign w1294 = w1169 & ~w1230;
assign w1295 = ~w1199 & w1293;
assign w1296 = w1294 & w1295;
assign w1297 = w1106 & w1296;
assign w1298 = w1013 & w1297;
assign w1299 = ~pi057 & pi153;
assign w1300 = ~pi056 & pi152;
assign w1301 = ~w1299 & ~w1300;
assign w1302 = pi056 & ~pi152;
assign w1303 = pi055 & ~pi151;
assign w1304 = ~w1302 & ~w1303;
assign w1305 = ~w1301 & w1304;
assign w1306 = pi060 & ~pi156;
assign w1307 = pi061 & ~pi157;
assign w1308 = ~pi061 & pi157;
assign w1309 = pi062 & ~pi158;
assign w1310 = ~w1308 & w1309;
assign w1311 = ~w1306 & ~w1307;
assign w1312 = ~w1310 & w1311;
assign w1313 = ~pi060 & pi156;
assign w1314 = ~pi059 & pi155;
assign w1315 = ~pi058 & pi154;
assign w1316 = ~w1313 & ~w1314;
assign w1317 = ~w1315 & w1316;
assign w1318 = ~w1312 & w1317;
assign w1319 = pi057 & ~pi153;
assign w1320 = pi059 & ~pi155;
assign w1321 = pi058 & ~pi154;
assign w1322 = ~w1320 & ~w1321;
assign w1323 = ~w1315 & ~w1322;
assign w1324 = w1304 & ~w1319;
assign w1325 = ~w1323 & w1324;
assign w1326 = ~w1318 & w1325;
assign w1327 = ~w1305 & ~w1326;
assign w1328 = ~pi055 & pi151;
assign w1329 = w1327 & ~w1328;
assign w1330 = ~pi061 & pi165;
assign w1331 = pi062 & ~pi166;
assign w1332 = ~w1330 & w1331;
assign w1333 = pi061 & ~pi165;
assign w1334 = pi060 & ~pi164;
assign w1335 = ~w1333 & ~w1334;
assign w1336 = ~w1332 & w1335;
assign w1337 = ~pi060 & pi164;
assign w1338 = ~pi059 & pi163;
assign w1339 = ~w1337 & ~w1338;
assign w1340 = pi059 & ~pi163;
assign w1341 = pi058 & ~pi162;
assign w1342 = ~w1340 & ~w1341;
assign w1343 = (w1342 & w1336) | (w1342 & w16188) | (w1336 & w16188);
assign w1344 = ~pi058 & pi162;
assign w1345 = ~pi057 & pi161;
assign w1346 = ~w1344 & ~w1345;
assign w1347 = ~w1343 & w1346;
assign w1348 = pi055 & ~pi159;
assign w1349 = pi056 & ~pi160;
assign w1350 = pi057 & ~pi161;
assign w1351 = ~w1348 & ~w1349;
assign w1352 = ~w1350 & w1351;
assign w1353 = ~w1347 & w1352;
assign w1354 = ~pi055 & pi159;
assign w1355 = ~pi056 & pi160;
assign w1356 = ~w1348 & w1355;
assign w1357 = ~w1354 & ~w1356;
assign w1358 = ~w1353 & w1357;
assign w1359 = ~w1329 & ~w1358;
assign w1360 = ~pi055 & pi111;
assign w1361 = pi056 & ~pi112;
assign w1362 = pi055 & ~pi111;
assign w1363 = ~w1361 & ~w1362;
assign w1364 = ~w1360 & ~w1363;
assign w1365 = pi062 & ~pi118;
assign w1366 = pi061 & ~pi117;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = ~pi061 & pi117;
assign w1369 = ~pi060 & pi116;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = ~w1367 & w1370;
assign w1372 = pi060 & ~pi116;
assign w1373 = pi059 & ~pi115;
assign w1374 = ~w1372 & ~w1373;
assign w1375 = ~pi059 & pi115;
assign w1376 = ~pi058 & pi114;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = (w1377 & w1371) | (w1377 & w16189) | (w1371 & w16189);
assign w1379 = pi058 & ~pi114;
assign w1380 = pi057 & ~pi113;
assign w1381 = ~w1379 & ~w1380;
assign w1382 = ~w1378 & w1381;
assign w1383 = ~pi057 & pi113;
assign w1384 = ~pi056 & pi112;
assign w1385 = ~w1383 & ~w1384;
assign w1386 = ~w1360 & w1385;
assign w1387 = ~w1382 & w1386;
assign w1388 = ~w1364 & ~w1387;
assign w1389 = ~pi061 & pi109;
assign w1390 = pi062 & ~pi110;
assign w1391 = ~w1389 & w1390;
assign w1392 = pi061 & ~pi109;
assign w1393 = pi060 & ~pi108;
assign w1394 = ~w1392 & ~w1393;
assign w1395 = ~w1391 & w1394;
assign w1396 = ~pi060 & pi108;
assign w1397 = ~pi059 & pi107;
assign w1398 = ~w1396 & ~w1397;
assign w1399 = pi059 & ~pi107;
assign w1400 = pi058 & ~pi106;
assign w1401 = ~w1399 & ~w1400;
assign w1402 = (w1401 & w1395) | (w1401 & w16190) | (w1395 & w16190);
assign w1403 = ~pi058 & pi106;
assign w1404 = ~pi057 & pi105;
assign w1405 = ~w1403 & ~w1404;
assign w1406 = ~w1402 & w1405;
assign w1407 = pi055 & ~pi103;
assign w1408 = pi056 & ~pi104;
assign w1409 = pi057 & ~pi105;
assign w1410 = ~w1407 & ~w1408;
assign w1411 = ~w1409 & w1410;
assign w1412 = ~w1406 & w1411;
assign w1413 = ~pi055 & pi103;
assign w1414 = ~pi056 & pi104;
assign w1415 = ~w1407 & w1414;
assign w1416 = ~w1413 & ~w1415;
assign w1417 = ~w1412 & w1416;
assign w1418 = w1388 & ~w1417;
assign w1419 = w1359 & w1418;
assign w1420 = ~w950 & ~w951;
assign w1421 = w29 & ~w1420;
assign w1422 = w1419 & w1421;
assign w1423 = w1298 & w1422;
assign w1424 = ~pi055 & pi271;
assign w1425 = pi058 & ~pi274;
assign w1426 = pi057 & ~pi273;
assign w1427 = ~w1425 & ~w1426;
assign w1428 = ~pi057 & pi273;
assign w1429 = ~pi056 & pi272;
assign w1430 = ~w1428 & ~w1429;
assign w1431 = ~w1427 & w1430;
assign w1432 = pi062 & ~pi278;
assign w1433 = pi061 & ~pi277;
assign w1434 = ~w1432 & ~w1433;
assign w1435 = ~pi061 & pi277;
assign w1436 = ~pi060 & pi276;
assign w1437 = ~w1435 & ~w1436;
assign w1438 = ~w1434 & w1437;
assign w1439 = pi060 & ~pi276;
assign w1440 = pi059 & ~pi275;
assign w1441 = ~w1439 & ~w1440;
assign w1442 = ~w1438 & w1441;
assign w1443 = ~pi058 & pi274;
assign w1444 = ~pi059 & pi275;
assign w1445 = ~w1443 & ~w1444;
assign w1446 = w1430 & w1445;
assign w1447 = (~w1431 & w1442) | (~w1431 & w16191) | (w1442 & w16191);
assign w1448 = pi056 & ~pi272;
assign w1449 = pi055 & ~pi271;
assign w1450 = ~w1448 & ~w1449;
assign w1451 = w1447 & w1450;
assign w1452 = (~w1424 & ~w1447) | (~w1424 & w16991) | (~w1447 & w16991);
assign w1453 = ~pi055 & pi263;
assign w1454 = pi060 & ~pi268;
assign w1455 = pi061 & ~pi269;
assign w1456 = ~pi061 & pi269;
assign w1457 = pi062 & ~pi270;
assign w1458 = ~w1456 & w1457;
assign w1459 = ~w1454 & ~w1455;
assign w1460 = ~w1458 & w1459;
assign w1461 = ~pi059 & pi267;
assign w1462 = ~pi058 & pi266;
assign w1463 = ~pi057 & pi265;
assign w1464 = ~w1462 & ~w1463;
assign w1465 = ~pi060 & pi268;
assign w1466 = ~w1461 & ~w1465;
assign w1467 = w1464 & w1466;
assign w1468 = ~w1460 & w1467;
assign w1469 = pi056 & ~pi264;
assign w1470 = pi059 & ~pi267;
assign w1471 = pi058 & ~pi266;
assign w1472 = ~w1470 & ~w1471;
assign w1473 = w1464 & ~w1472;
assign w1474 = pi055 & ~pi263;
assign w1475 = pi057 & ~pi265;
assign w1476 = ~w1469 & ~w1474;
assign w1477 = ~w1475 & w1476;
assign w1478 = ~w1473 & w1477;
assign w1479 = ~w1468 & w1478;
assign w1480 = ~pi056 & pi264;
assign w1481 = ~w1474 & w1480;
assign w1482 = ~w1479 & ~w1481;
assign w1483 = ~w1479 & w16992;
assign w1484 = ~w1452 & ~w1483;
assign w1485 = ~pi057 & pi249;
assign w1486 = ~pi056 & pi248;
assign w1487 = ~w1485 & ~w1486;
assign w1488 = pi056 & ~pi248;
assign w1489 = pi055 & ~pi247;
assign w1490 = ~w1488 & ~w1489;
assign w1491 = ~w1487 & w1490;
assign w1492 = pi060 & ~pi252;
assign w1493 = pi061 & ~pi253;
assign w1494 = ~pi061 & pi253;
assign w1495 = pi062 & ~pi254;
assign w1496 = ~w1494 & w1495;
assign w1497 = ~w1492 & ~w1493;
assign w1498 = ~w1496 & w1497;
assign w1499 = ~pi060 & pi252;
assign w1500 = ~pi059 & pi251;
assign w1501 = ~pi058 & pi250;
assign w1502 = ~w1499 & ~w1500;
assign w1503 = ~w1501 & w1502;
assign w1504 = ~w1498 & w1503;
assign w1505 = pi057 & ~pi249;
assign w1506 = pi059 & ~pi251;
assign w1507 = pi058 & ~pi250;
assign w1508 = ~w1506 & ~w1507;
assign w1509 = ~w1501 & ~w1508;
assign w1510 = w1490 & ~w1505;
assign w1511 = ~w1509 & w1510;
assign w1512 = ~w1504 & w1511;
assign w1513 = ~w1491 & ~w1512;
assign w1514 = ~pi055 & pi247;
assign w1515 = ~w1512 & w16993;
assign w1516 = ~pi055 & pi255;
assign w1517 = pi060 & ~pi260;
assign w1518 = pi061 & ~pi261;
assign w1519 = ~pi061 & pi261;
assign w1520 = pi062 & ~pi262;
assign w1521 = ~w1519 & w1520;
assign w1522 = ~w1517 & ~w1518;
assign w1523 = ~w1521 & w1522;
assign w1524 = ~pi059 & pi259;
assign w1525 = ~pi058 & pi258;
assign w1526 = ~pi057 & pi257;
assign w1527 = ~w1525 & ~w1526;
assign w1528 = ~pi060 & pi260;
assign w1529 = ~w1524 & ~w1528;
assign w1530 = w1527 & w1529;
assign w1531 = ~w1523 & w1530;
assign w1532 = pi057 & ~pi257;
assign w1533 = pi059 & ~pi259;
assign w1534 = pi058 & ~pi258;
assign w1535 = ~w1533 & ~w1534;
assign w1536 = w1527 & ~w1535;
assign w1537 = pi055 & ~pi255;
assign w1538 = pi056 & ~pi256;
assign w1539 = ~w1532 & ~w1537;
assign w1540 = ~w1538 & w1539;
assign w1541 = ~w1536 & w1540;
assign w1542 = ~w1531 & w1541;
assign w1543 = ~pi056 & pi256;
assign w1544 = ~w1537 & w1543;
assign w1545 = ~w1542 & ~w1544;
assign w1546 = ~w1542 & w16994;
assign w1547 = ~w1515 & ~w1546;
assign w1548 = w1484 & w1547;
assign w1549 = pi061 & ~pi237;
assign w1550 = pi060 & ~pi236;
assign w1551 = ~pi061 & pi237;
assign w1552 = pi062 & ~pi238;
assign w1553 = ~w1551 & w1552;
assign w1554 = ~w1549 & ~w1550;
assign w1555 = ~w1553 & w1554;
assign w1556 = ~pi059 & pi235;
assign w1557 = ~pi058 & pi234;
assign w1558 = ~pi057 & pi233;
assign w1559 = ~w1557 & ~w1558;
assign w1560 = ~pi060 & pi236;
assign w1561 = ~w1556 & ~w1560;
assign w1562 = w1559 & w1561;
assign w1563 = ~w1555 & w1562;
assign w1564 = pi055 & ~pi231;
assign w1565 = pi059 & ~pi235;
assign w1566 = pi058 & ~pi234;
assign w1567 = ~w1565 & ~w1566;
assign w1568 = w1559 & ~w1567;
assign w1569 = pi056 & ~pi232;
assign w1570 = pi057 & ~pi233;
assign w1571 = ~w1564 & ~w1569;
assign w1572 = ~w1570 & w1571;
assign w1573 = ~w1568 & w1572;
assign w1574 = ~w1563 & w1573;
assign w1575 = ~pi055 & pi231;
assign w1576 = ~pi056 & pi232;
assign w1577 = ~w1564 & w1576;
assign w1578 = ~w1575 & ~w1577;
assign w1579 = ~w1574 & w1578;
assign w1580 = ~pi055 & pi239;
assign w1581 = ~pi061 & pi245;
assign w1582 = pi062 & ~pi246;
assign w1583 = ~w1581 & w1582;
assign w1584 = pi061 & ~pi245;
assign w1585 = pi060 & ~pi244;
assign w1586 = ~w1584 & ~w1585;
assign w1587 = ~w1583 & w1586;
assign w1588 = ~pi058 & pi242;
assign w1589 = ~pi057 & pi241;
assign w1590 = ~w1588 & ~w1589;
assign w1591 = ~pi060 & pi244;
assign w1592 = ~pi059 & pi243;
assign w1593 = ~w1591 & ~w1592;
assign w1594 = w1590 & w1593;
assign w1595 = ~w1587 & w1594;
assign w1596 = pi059 & ~pi243;
assign w1597 = pi058 & ~pi242;
assign w1598 = ~w1596 & ~w1597;
assign w1599 = w1590 & ~w1598;
assign w1600 = pi057 & ~pi241;
assign w1601 = pi055 & ~pi239;
assign w1602 = pi056 & ~pi240;
assign w1603 = ~w1600 & ~w1601;
assign w1604 = ~w1602 & w1603;
assign w1605 = ~w1599 & w1604;
assign w1606 = ~w1595 & w1605;
assign w1607 = ~pi056 & pi240;
assign w1608 = ~w1601 & w1607;
assign w1609 = ~w1606 & ~w1608;
assign w1610 = ~w1606 & w16192;
assign w1611 = ~w1579 & ~w1610;
assign w1612 = ~pi055 & pi215;
assign w1613 = pi056 & ~pi216;
assign w1614 = pi055 & ~pi215;
assign w1615 = ~w1613 & ~w1614;
assign w1616 = ~w1612 & ~w1615;
assign w1617 = pi062 & ~pi222;
assign w1618 = pi061 & ~pi221;
assign w1619 = ~w1617 & ~w1618;
assign w1620 = ~pi061 & pi221;
assign w1621 = ~pi060 & pi220;
assign w1622 = ~w1620 & ~w1621;
assign w1623 = ~w1619 & w1622;
assign w1624 = pi060 & ~pi220;
assign w1625 = pi059 & ~pi219;
assign w1626 = ~w1624 & ~w1625;
assign w1627 = ~pi059 & pi219;
assign w1628 = ~pi058 & pi218;
assign w1629 = ~w1627 & ~w1628;
assign w1630 = (w1629 & w1623) | (w1629 & w16193) | (w1623 & w16193);
assign w1631 = pi058 & ~pi218;
assign w1632 = pi057 & ~pi217;
assign w1633 = ~w1631 & ~w1632;
assign w1634 = ~w1630 & w1633;
assign w1635 = ~pi057 & pi217;
assign w1636 = ~pi056 & pi216;
assign w1637 = ~w1635 & ~w1636;
assign w1638 = ~w1612 & w1637;
assign w1639 = (w1638 & w1630) | (w1638 & w16995) | (w1630 & w16995);
assign w1640 = ~w1616 & ~w1639;
assign w1641 = w1611 & w1640;
assign w1642 = pi055 & ~pi183;
assign w1643 = ~pi061 & pi189;
assign w1644 = pi062 & ~pi190;
assign w1645 = ~w1643 & w1644;
assign w1646 = pi061 & ~pi189;
assign w1647 = pi060 & ~pi188;
assign w1648 = ~w1646 & ~w1647;
assign w1649 = ~w1645 & w1648;
assign w1650 = ~pi060 & pi188;
assign w1651 = ~pi059 & pi187;
assign w1652 = ~w1650 & ~w1651;
assign w1653 = pi059 & ~pi187;
assign w1654 = pi058 & ~pi186;
assign w1655 = ~w1653 & ~w1654;
assign w1656 = (w1655 & w1649) | (w1655 & w16194) | (w1649 & w16194);
assign w1657 = ~pi058 & pi186;
assign w1658 = ~pi057 & pi185;
assign w1659 = ~w1657 & ~w1658;
assign w1660 = pi057 & ~pi185;
assign w1661 = pi056 & ~pi184;
assign w1662 = ~w1660 & ~w1661;
assign w1663 = (w1662 & w1656) | (w1662 & w16996) | (w1656 & w16996);
assign w1664 = ~pi056 & pi184;
assign w1665 = ~pi055 & pi183;
assign w1666 = ~w1664 & ~w1665;
assign w1667 = ~w1663 & w1666;
assign w1668 = ~w1642 & ~w1667;
assign w1669 = w1641 & w1668;
assign w1670 = w1548 & w1669;
assign w1671 = ~pi055 & pi223;
assign w1672 = pi056 & ~pi224;
assign w1673 = pi055 & ~pi223;
assign w1674 = ~w1672 & ~w1673;
assign w1675 = ~w1671 & ~w1674;
assign w1676 = pi062 & ~pi230;
assign w1677 = pi061 & ~pi229;
assign w1678 = ~w1676 & ~w1677;
assign w1679 = ~pi061 & pi229;
assign w1680 = ~pi060 & pi228;
assign w1681 = ~w1679 & ~w1680;
assign w1682 = ~w1678 & w1681;
assign w1683 = pi060 & ~pi228;
assign w1684 = pi059 & ~pi227;
assign w1685 = ~w1683 & ~w1684;
assign w1686 = ~pi059 & pi227;
assign w1687 = ~pi058 & pi226;
assign w1688 = ~w1686 & ~w1687;
assign w1689 = (w1688 & w1682) | (w1688 & w16195) | (w1682 & w16195);
assign w1690 = pi058 & ~pi226;
assign w1691 = pi057 & ~pi225;
assign w1692 = ~w1690 & ~w1691;
assign w1693 = ~w1689 & w1692;
assign w1694 = ~pi057 & pi225;
assign w1695 = ~pi056 & pi224;
assign w1696 = ~w1694 & ~w1695;
assign w1697 = ~w1671 & w1696;
assign w1698 = (w1697 & w1689) | (w1697 & w16997) | (w1689 & w16997);
assign w1699 = ~w1675 & ~w1698;
assign w1700 = pi062 & ~pi206;
assign w1701 = pi061 & ~pi205;
assign w1702 = ~w1700 & ~w1701;
assign w1703 = ~pi061 & pi205;
assign w1704 = ~pi060 & pi204;
assign w1705 = ~w1703 & ~w1704;
assign w1706 = ~w1702 & w1705;
assign w1707 = pi060 & ~pi204;
assign w1708 = pi059 & ~pi203;
assign w1709 = ~w1707 & ~w1708;
assign w1710 = ~pi059 & pi203;
assign w1711 = ~pi058 & pi202;
assign w1712 = ~w1710 & ~w1711;
assign w1713 = (w1712 & w1706) | (w1712 & w16196) | (w1706 & w16196);
assign w1714 = pi058 & ~pi202;
assign w1715 = pi057 & ~pi201;
assign w1716 = ~w1714 & ~w1715;
assign w1717 = ~pi055 & pi199;
assign w1718 = ~pi056 & pi200;
assign w1719 = ~pi057 & pi201;
assign w1720 = ~w1717 & ~w1718;
assign w1721 = ~w1719 & w1720;
assign w1722 = (w1721 & w1713) | (w1721 & w16998) | (w1713 & w16998);
assign w1723 = pi055 & ~pi199;
assign w1724 = pi056 & ~pi200;
assign w1725 = ~w1717 & w1724;
assign w1726 = ~w1723 & ~w1725;
assign w1727 = ~w1722 & w1726;
assign w1728 = w1699 & w1727;
assign w1729 = ~pi055 & pi207;
assign w1730 = pi062 & ~pi214;
assign w1731 = pi061 & ~pi213;
assign w1732 = ~w1730 & ~w1731;
assign w1733 = ~pi061 & pi213;
assign w1734 = ~pi060 & pi212;
assign w1735 = ~w1733 & ~w1734;
assign w1736 = ~w1732 & w1735;
assign w1737 = pi060 & ~pi212;
assign w1738 = pi059 & ~pi211;
assign w1739 = ~w1737 & ~w1738;
assign w1740 = ~pi059 & pi211;
assign w1741 = ~pi058 & pi210;
assign w1742 = ~w1740 & ~w1741;
assign w1743 = (w1742 & w1736) | (w1742 & w16197) | (w1736 & w16197);
assign w1744 = pi058 & ~pi210;
assign w1745 = pi057 & ~pi209;
assign w1746 = ~w1744 & ~w1745;
assign w1747 = ~pi057 & pi209;
assign w1748 = ~pi056 & pi208;
assign w1749 = ~w1747 & ~w1748;
assign w1750 = (w1749 & w1743) | (w1749 & w16999) | (w1743 & w16999);
assign w1751 = pi056 & ~pi208;
assign w1752 = pi055 & ~pi207;
assign w1753 = ~w1751 & ~w1752;
assign w1754 = ~w1750 & w1753;
assign w1755 = ~w1729 & ~w1754;
assign w1756 = w1728 & ~w1755;
assign w1757 = w467 & w1756;
assign w1758 = w1670 & w1757;
assign w1759 = w1423 & w1758;
assign w1760 = pi003 & w1759;
assign w1761 = ~pi002 & ~w29;
assign w1762 = ~pi001 & w29;
assign w1763 = ~w1761 & ~w1762;
assign w1764 = w918 & w1763;
assign w1765 = ~w956 & ~w1764;
assign w1766 = ~w1760 & w1765;
assign w1767 = ~w404 & ~w918;
assign w1768 = ~pi071 & pi239;
assign w1769 = pi072 & ~pi240;
assign w1770 = pi071 & ~pi239;
assign w1771 = ~w1769 & ~w1770;
assign w1772 = ~w1768 & ~w1771;
assign w1773 = pi078 & ~pi246;
assign w1774 = pi077 & ~pi245;
assign w1775 = ~w1773 & ~w1774;
assign w1776 = ~pi077 & pi245;
assign w1777 = ~pi076 & pi244;
assign w1778 = ~w1776 & ~w1777;
assign w1779 = ~w1775 & w1778;
assign w1780 = pi076 & ~pi244;
assign w1781 = pi075 & ~pi243;
assign w1782 = ~w1780 & ~w1781;
assign w1783 = ~pi075 & pi243;
assign w1784 = ~pi074 & pi242;
assign w1785 = ~w1783 & ~w1784;
assign w1786 = (w1785 & w1779) | (w1785 & w16198) | (w1779 & w16198);
assign w1787 = pi074 & ~pi242;
assign w1788 = pi073 & ~pi241;
assign w1789 = ~w1787 & ~w1788;
assign w1790 = ~w1786 & w1789;
assign w1791 = ~pi073 & pi241;
assign w1792 = ~pi072 & pi240;
assign w1793 = ~w1791 & ~w1792;
assign w1794 = ~w1768 & w1793;
assign w1795 = ~w1790 & w1794;
assign w1796 = ~w1772 & ~w1795;
assign w1797 = ~pi071 & pi231;
assign w1798 = pi072 & ~pi232;
assign w1799 = pi071 & ~pi231;
assign w1800 = ~w1798 & ~w1799;
assign w1801 = ~w1797 & ~w1800;
assign w1802 = pi078 & ~pi238;
assign w1803 = pi077 & ~pi237;
assign w1804 = ~w1802 & ~w1803;
assign w1805 = ~pi077 & pi237;
assign w1806 = ~pi076 & pi236;
assign w1807 = ~w1805 & ~w1806;
assign w1808 = ~w1804 & w1807;
assign w1809 = pi076 & ~pi236;
assign w1810 = pi075 & ~pi235;
assign w1811 = ~w1809 & ~w1810;
assign w1812 = ~pi075 & pi235;
assign w1813 = ~pi074 & pi234;
assign w1814 = ~w1812 & ~w1813;
assign w1815 = (w1814 & w1808) | (w1814 & w16199) | (w1808 & w16199);
assign w1816 = pi074 & ~pi234;
assign w1817 = pi073 & ~pi233;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = ~w1815 & w1818;
assign w1820 = ~pi073 & pi233;
assign w1821 = ~pi072 & pi232;
assign w1822 = ~w1820 & ~w1821;
assign w1823 = ~w1797 & w1822;
assign w1824 = ~w1819 & w1823;
assign w1825 = ~w1801 & ~w1824;
assign w1826 = w1796 & w1825;
assign w1827 = pi072 & ~pi264;
assign w1828 = pi071 & ~pi263;
assign w1829 = ~w1827 & ~w1828;
assign w1830 = ~pi071 & pi263;
assign w1831 = ~w1829 & ~w1830;
assign w1832 = pi078 & ~pi270;
assign w1833 = pi077 & ~pi269;
assign w1834 = ~w1832 & ~w1833;
assign w1835 = ~pi077 & pi269;
assign w1836 = ~pi076 & pi268;
assign w1837 = ~w1835 & ~w1836;
assign w1838 = ~w1834 & w1837;
assign w1839 = pi076 & ~pi268;
assign w1840 = pi075 & ~pi267;
assign w1841 = ~w1839 & ~w1840;
assign w1842 = ~pi075 & pi267;
assign w1843 = ~pi074 & pi266;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = (w1844 & w1838) | (w1844 & w16200) | (w1838 & w16200);
assign w1846 = pi074 & ~pi266;
assign w1847 = pi073 & ~pi265;
assign w1848 = ~w1846 & ~w1847;
assign w1849 = ~w1845 & w1848;
assign w1850 = ~pi073 & pi265;
assign w1851 = ~pi072 & pi264;
assign w1852 = ~w1850 & ~w1851;
assign w1853 = ~w1830 & w1852;
assign w1854 = ~w1849 & w1853;
assign w1855 = ~w1831 & ~w1854;
assign w1856 = pi074 & ~pi250;
assign w1857 = ~pi075 & pi251;
assign w1858 = ~pi074 & pi250;
assign w1859 = ~w1857 & ~w1858;
assign w1860 = pi076 & ~pi252;
assign w1861 = pi075 & ~pi251;
assign w1862 = ~w1860 & ~w1861;
assign w1863 = w1859 & ~w1862;
assign w1864 = pi072 & ~pi248;
assign w1865 = pi071 & ~pi247;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = pi073 & ~pi249;
assign w1868 = ~pi077 & pi253;
assign w1869 = pi077 & ~pi253;
assign w1870 = pi078 & ~pi254;
assign w1871 = ~w1869 & ~w1870;
assign w1872 = ~pi076 & pi252;
assign w1873 = ~w1868 & ~w1872;
assign w1874 = w1859 & w1873;
assign w1875 = ~w1871 & w1874;
assign w1876 = ~w1856 & ~w1867;
assign w1877 = w1866 & w1876;
assign w1878 = ~w1863 & w1877;
assign w1879 = ~w1875 & w1878;
assign w1880 = ~pi071 & pi247;
assign w1881 = ~pi073 & pi249;
assign w1882 = ~pi072 & pi248;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = w1866 & ~w1883;
assign w1885 = ~w1880 & ~w1884;
assign w1886 = ~w1879 & w1885;
assign w1887 = ~pi075 & pi259;
assign w1888 = ~pi074 & pi258;
assign w1889 = ~w1887 & ~w1888;
assign w1890 = pi076 & ~pi260;
assign w1891 = pi075 & ~pi259;
assign w1892 = ~w1890 & ~w1891;
assign w1893 = w1889 & ~w1892;
assign w1894 = pi072 & ~pi256;
assign w1895 = pi071 & ~pi255;
assign w1896 = ~w1894 & ~w1895;
assign w1897 = pi074 & ~pi258;
assign w1898 = pi073 & ~pi257;
assign w1899 = pi078 & ~pi262;
assign w1900 = pi077 & ~pi261;
assign w1901 = ~w1899 & ~w1900;
assign w1902 = ~pi077 & pi261;
assign w1903 = ~pi076 & pi260;
assign w1904 = ~w1902 & ~w1903;
assign w1905 = w1889 & w1904;
assign w1906 = ~w1901 & w1905;
assign w1907 = ~w1897 & ~w1898;
assign w1908 = w1896 & w1907;
assign w1909 = ~w1893 & w1908;
assign w1910 = ~w1906 & w1909;
assign w1911 = ~pi073 & pi257;
assign w1912 = ~pi072 & pi256;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = w1896 & ~w1913;
assign w1915 = ~w1910 & ~w1914;
assign w1916 = ~pi071 & pi255;
assign w1917 = ~w1910 & w16201;
assign w1918 = ~w1886 & ~w1917;
assign w1919 = w1855 & w1918;
assign w1920 = w1826 & w1919;
assign w1921 = ~pi071 & pi135;
assign w1922 = pi075 & ~pi139;
assign w1923 = pi076 & ~pi140;
assign w1924 = ~pi076 & pi140;
assign w1925 = pi078 & ~pi142;
assign w1926 = pi077 & ~pi141;
assign w1927 = ~w1925 & ~w1926;
assign w1928 = ~pi077 & pi141;
assign w1929 = ~w1924 & ~w1928;
assign w1930 = ~w1927 & w1929;
assign w1931 = ~w1922 & ~w1923;
assign w1932 = ~w1930 & w1931;
assign w1933 = ~pi075 & pi139;
assign w1934 = ~pi074 & pi138;
assign w1935 = ~w1933 & ~w1934;
assign w1936 = ~w1932 & w1935;
assign w1937 = pi074 & ~pi138;
assign w1938 = pi073 & ~pi137;
assign w1939 = ~w1937 & ~w1938;
assign w1940 = ~w1936 & w1939;
assign w1941 = ~pi073 & pi137;
assign w1942 = ~pi072 & pi136;
assign w1943 = ~w1941 & ~w1942;
assign w1944 = ~w1940 & w1943;
assign w1945 = pi072 & ~pi136;
assign w1946 = pi071 & ~pi135;
assign w1947 = ~w1945 & ~w1946;
assign w1948 = ~w1944 & w1947;
assign w1949 = ~w1921 & ~w1948;
assign w1950 = w1920 & ~w1949;
assign w1951 = ~pi075 & pi211;
assign w1952 = ~pi074 & pi210;
assign w1953 = ~w1951 & ~w1952;
assign w1954 = pi076 & ~pi212;
assign w1955 = pi075 & ~pi211;
assign w1956 = ~w1954 & ~w1955;
assign w1957 = w1953 & ~w1956;
assign w1958 = pi072 & ~pi208;
assign w1959 = pi071 & ~pi207;
assign w1960 = ~w1958 & ~w1959;
assign w1961 = pi074 & ~pi210;
assign w1962 = pi073 & ~pi209;
assign w1963 = pi078 & ~pi214;
assign w1964 = pi077 & ~pi213;
assign w1965 = ~w1963 & ~w1964;
assign w1966 = ~pi077 & pi213;
assign w1967 = ~pi076 & pi212;
assign w1968 = ~w1966 & ~w1967;
assign w1969 = w1953 & w1968;
assign w1970 = ~w1965 & w1969;
assign w1971 = ~w1961 & ~w1962;
assign w1972 = w1960 & w1971;
assign w1973 = ~w1957 & w1972;
assign w1974 = ~w1970 & w1973;
assign w1975 = ~pi073 & pi209;
assign w1976 = ~pi072 & pi208;
assign w1977 = ~w1975 & ~w1976;
assign w1978 = w1960 & ~w1977;
assign w1979 = ~w1974 & ~w1978;
assign w1980 = ~pi071 & pi207;
assign w1981 = ~w1974 & w16202;
assign w1982 = pi078 & ~pi206;
assign w1983 = pi077 & ~pi205;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = ~pi077 & pi205;
assign w1986 = ~pi076 & pi204;
assign w1987 = ~w1985 & ~w1986;
assign w1988 = ~w1984 & w1987;
assign w1989 = pi074 & ~pi202;
assign w1990 = pi073 & ~pi201;
assign w1991 = ~w1989 & ~w1990;
assign w1992 = pi076 & ~pi204;
assign w1993 = pi075 & ~pi203;
assign w1994 = ~w1992 & ~w1993;
assign w1995 = w1991 & w1994;
assign w1996 = ~w1988 & w1995;
assign w1997 = ~pi075 & pi203;
assign w1998 = ~pi074 & pi202;
assign w1999 = ~w1997 & ~w1998;
assign w2000 = w1991 & ~w1999;
assign w2001 = ~pi073 & pi201;
assign w2002 = ~pi072 & pi200;
assign w2003 = ~w2001 & ~w2002;
assign w2004 = ~w2000 & w2003;
assign w2005 = ~w1996 & w2004;
assign w2006 = pi072 & ~pi200;
assign w2007 = pi071 & ~pi199;
assign w2008 = ~w2006 & ~w2007;
assign w2009 = ~w2005 & w2008;
assign w2010 = ~pi071 & pi199;
assign w2011 = (~w2010 & w2005) | (~w2010 & w16203) | (w2005 & w16203);
assign w2012 = ~w1981 & ~w2011;
assign w2013 = ~pi076 & pi188;
assign w2014 = pi078 & ~pi190;
assign w2015 = pi077 & ~pi189;
assign w2016 = ~w2014 & ~w2015;
assign w2017 = ~pi077 & pi189;
assign w2018 = ~w2013 & ~w2017;
assign w2019 = ~w2016 & w2018;
assign w2020 = pi076 & ~pi188;
assign w2021 = pi074 & ~pi186;
assign w2022 = pi073 & ~pi185;
assign w2023 = ~w2021 & ~w2022;
assign w2024 = pi075 & ~pi187;
assign w2025 = ~w2020 & ~w2024;
assign w2026 = w2023 & w2025;
assign w2027 = ~w2019 & w2026;
assign w2028 = ~pi073 & pi185;
assign w2029 = ~pi075 & pi187;
assign w2030 = ~pi074 & pi186;
assign w2031 = ~w2029 & ~w2030;
assign w2032 = w2023 & ~w2031;
assign w2033 = ~pi072 & pi184;
assign w2034 = ~w2028 & ~w2033;
assign w2035 = ~w2032 & w2034;
assign w2036 = ~w2027 & w2035;
assign w2037 = pi072 & ~pi184;
assign w2038 = pi071 & ~pi183;
assign w2039 = ~w2037 & ~w2038;
assign w2040 = ~w2036 & w2039;
assign w2041 = ~pi071 & pi183;
assign w2042 = ~w2040 & ~w2041;
assign w2043 = w2012 & ~w2042;
assign w2044 = pi078 & ~pi222;
assign w2045 = pi077 & ~pi221;
assign w2046 = ~w2044 & ~w2045;
assign w2047 = ~pi077 & pi221;
assign w2048 = ~pi076 & pi220;
assign w2049 = ~w2047 & ~w2048;
assign w2050 = ~w2046 & w2049;
assign w2051 = pi074 & ~pi218;
assign w2052 = pi073 & ~pi217;
assign w2053 = ~w2051 & ~w2052;
assign w2054 = pi076 & ~pi220;
assign w2055 = pi075 & ~pi219;
assign w2056 = ~w2054 & ~w2055;
assign w2057 = w2053 & w2056;
assign w2058 = ~w2050 & w2057;
assign w2059 = ~pi075 & pi219;
assign w2060 = ~pi074 & pi218;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = w2053 & ~w2061;
assign w2063 = ~pi073 & pi217;
assign w2064 = ~pi072 & pi216;
assign w2065 = ~w2063 & ~w2064;
assign w2066 = ~w2062 & w2065;
assign w2067 = ~w2058 & w2066;
assign w2068 = pi072 & ~pi216;
assign w2069 = pi071 & ~pi215;
assign w2070 = ~w2068 & ~w2069;
assign w2071 = ~w2067 & w2070;
assign w2072 = ~pi071 & pi215;
assign w2073 = (~w2072 & w2067) | (~w2072 & w16204) | (w2067 & w16204);
assign w2074 = pi078 & ~pi278;
assign w2075 = pi077 & ~pi277;
assign w2076 = ~w2074 & ~w2075;
assign w2077 = ~pi077 & pi277;
assign w2078 = ~pi076 & pi276;
assign w2079 = ~w2077 & ~w2078;
assign w2080 = ~w2076 & w2079;
assign w2081 = pi074 & ~pi274;
assign w2082 = pi073 & ~pi273;
assign w2083 = ~w2081 & ~w2082;
assign w2084 = pi076 & ~pi276;
assign w2085 = pi075 & ~pi275;
assign w2086 = ~w2084 & ~w2085;
assign w2087 = w2083 & w2086;
assign w2088 = ~w2080 & w2087;
assign w2089 = ~pi075 & pi275;
assign w2090 = ~pi074 & pi274;
assign w2091 = ~w2089 & ~w2090;
assign w2092 = w2083 & ~w2091;
assign w2093 = ~pi073 & pi273;
assign w2094 = ~pi072 & pi272;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = ~w2092 & w2095;
assign w2097 = ~w2088 & w2096;
assign w2098 = pi072 & ~pi272;
assign w2099 = pi071 & ~pi271;
assign w2100 = ~w2098 & ~w2099;
assign w2101 = ~w2097 & w2100;
assign w2102 = ~pi071 & pi271;
assign w2103 = (~w2102 & w2097) | (~w2102 & w16205) | (w2097 & w16205);
assign w2104 = ~w2073 & ~w2103;
assign w2105 = pi078 & ~pi174;
assign w2106 = pi077 & ~pi173;
assign w2107 = ~w2105 & ~w2106;
assign w2108 = ~pi077 & pi173;
assign w2109 = ~pi076 & pi172;
assign w2110 = ~w2108 & ~w2109;
assign w2111 = ~w2107 & w2110;
assign w2112 = pi074 & ~pi170;
assign w2113 = pi073 & ~pi169;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = pi076 & ~pi172;
assign w2116 = pi075 & ~pi171;
assign w2117 = ~w2115 & ~w2116;
assign w2118 = w2114 & w2117;
assign w2119 = ~w2111 & w2118;
assign w2120 = ~pi075 & pi171;
assign w2121 = ~pi074 & pi170;
assign w2122 = ~w2120 & ~w2121;
assign w2123 = w2114 & ~w2122;
assign w2124 = ~pi073 & pi169;
assign w2125 = ~pi072 & pi168;
assign w2126 = ~w2124 & ~w2125;
assign w2127 = ~w2123 & w2126;
assign w2128 = ~w2119 & w2127;
assign w2129 = pi072 & ~pi168;
assign w2130 = pi071 & ~pi167;
assign w2131 = ~w2129 & ~w2130;
assign w2132 = ~w2128 & w2131;
assign w2133 = ~pi071 & pi167;
assign w2134 = (~w2133 & w2128) | (~w2133 & w16206) | (w2128 & w16206);
assign w2135 = pi078 & ~pi158;
assign w2136 = pi077 & ~pi157;
assign w2137 = ~w2135 & ~w2136;
assign w2138 = ~pi077 & pi157;
assign w2139 = ~pi076 & pi156;
assign w2140 = ~w2138 & ~w2139;
assign w2141 = ~w2137 & w2140;
assign w2142 = pi074 & ~pi154;
assign w2143 = pi073 & ~pi153;
assign w2144 = ~w2142 & ~w2143;
assign w2145 = pi076 & ~pi156;
assign w2146 = pi075 & ~pi155;
assign w2147 = ~w2145 & ~w2146;
assign w2148 = w2144 & w2147;
assign w2149 = ~w2141 & w2148;
assign w2150 = ~pi075 & pi155;
assign w2151 = ~pi074 & pi154;
assign w2152 = ~w2150 & ~w2151;
assign w2153 = w2144 & ~w2152;
assign w2154 = ~pi073 & pi153;
assign w2155 = ~pi072 & pi152;
assign w2156 = ~w2154 & ~w2155;
assign w2157 = ~w2153 & w2156;
assign w2158 = ~w2149 & w2157;
assign w2159 = pi072 & ~pi152;
assign w2160 = pi071 & ~pi151;
assign w2161 = ~w2159 & ~w2160;
assign w2162 = ~w2158 & w2161;
assign w2163 = ~pi071 & pi151;
assign w2164 = (~w2163 & w2158) | (~w2163 & w16207) | (w2158 & w16207);
assign w2165 = ~w2134 & ~w2164;
assign w2166 = w2104 & w2165;
assign w2167 = w2043 & w2166;
assign w2168 = ~pi071 & pi223;
assign w2169 = ~pi075 & pi227;
assign w2170 = ~pi074 & pi226;
assign w2171 = ~w2169 & ~w2170;
assign w2172 = pi076 & ~pi228;
assign w2173 = pi075 & ~pi227;
assign w2174 = ~w2172 & ~w2173;
assign w2175 = w2171 & ~w2174;
assign w2176 = pi071 & ~pi223;
assign w2177 = pi072 & ~pi224;
assign w2178 = ~w2176 & ~w2177;
assign w2179 = pi074 & ~pi226;
assign w2180 = pi073 & ~pi225;
assign w2181 = pi078 & ~pi230;
assign w2182 = pi077 & ~pi229;
assign w2183 = ~w2181 & ~w2182;
assign w2184 = ~pi077 & pi229;
assign w2185 = ~pi076 & pi228;
assign w2186 = ~w2184 & ~w2185;
assign w2187 = w2171 & w2186;
assign w2188 = ~w2183 & w2187;
assign w2189 = ~w2179 & ~w2180;
assign w2190 = w2178 & w2189;
assign w2191 = ~w2175 & w2190;
assign w2192 = ~w2188 & w2191;
assign w2193 = ~pi073 & pi225;
assign w2194 = ~pi072 & pi224;
assign w2195 = ~w2193 & ~w2194;
assign w2196 = w2178 & ~w2195;
assign w2197 = ~w2192 & ~w2196;
assign w2198 = ~w2192 & w16208;
assign w2199 = ~pi075 & pi131;
assign w2200 = ~pi074 & pi130;
assign w2201 = ~w2199 & ~w2200;
assign w2202 = pi074 & ~pi130;
assign w2203 = pi073 & ~pi129;
assign w2204 = ~w2202 & ~w2203;
assign w2205 = ~w2201 & w2204;
assign w2206 = pi078 & ~pi134;
assign w2207 = pi077 & ~pi133;
assign w2208 = ~w2206 & ~w2207;
assign w2209 = ~pi077 & pi133;
assign w2210 = ~pi076 & pi132;
assign w2211 = ~w2209 & ~w2210;
assign w2212 = ~w2208 & w2211;
assign w2213 = pi076 & ~pi132;
assign w2214 = pi075 & ~pi131;
assign w2215 = ~w2213 & ~w2214;
assign w2216 = w2204 & w2215;
assign w2217 = ~w2212 & w2216;
assign w2218 = ~w2205 & ~w2217;
assign w2219 = ~pi071 & pi127;
assign w2220 = ~pi073 & pi129;
assign w2221 = ~pi072 & pi128;
assign w2222 = ~w2220 & ~w2221;
assign w2223 = ~w2219 & w2222;
assign w2224 = ~w2217 & w16209;
assign w2225 = pi072 & ~pi128;
assign w2226 = pi071 & ~pi127;
assign w2227 = ~w2225 & ~w2226;
assign w2228 = ~w2219 & ~w2227;
assign w2229 = ~w2224 & ~w2228;
assign w2230 = ~w2198 & w2229;
assign w2231 = ~pi071 & pi111;
assign w2232 = pi078 & ~pi118;
assign w2233 = pi077 & ~pi117;
assign w2234 = ~w2232 & ~w2233;
assign w2235 = ~pi076 & pi116;
assign w2236 = ~pi077 & pi117;
assign w2237 = ~w2235 & ~w2236;
assign w2238 = ~w2234 & w2237;
assign w2239 = pi074 & ~pi114;
assign w2240 = pi073 & ~pi113;
assign w2241 = ~w2239 & ~w2240;
assign w2242 = pi076 & ~pi116;
assign w2243 = pi075 & ~pi115;
assign w2244 = ~w2242 & ~w2243;
assign w2245 = w2241 & w2244;
assign w2246 = ~w2238 & w2245;
assign w2247 = ~pi075 & pi115;
assign w2248 = ~pi074 & pi114;
assign w2249 = ~w2247 & ~w2248;
assign w2250 = w2241 & ~w2249;
assign w2251 = ~pi073 & pi113;
assign w2252 = ~pi072 & pi112;
assign w2253 = ~w2251 & ~w2252;
assign w2254 = ~w2250 & w2253;
assign w2255 = ~w2246 & w2254;
assign w2256 = pi072 & ~pi112;
assign w2257 = pi071 & ~pi111;
assign w2258 = ~w2256 & ~w2257;
assign w2259 = ~w2255 & w2258;
assign w2260 = (~w2231 & w2255) | (~w2231 & w16210) | (w2255 & w16210);
assign w2261 = ~pi077 & pi149;
assign w2262 = pi078 & ~pi150;
assign w2263 = ~w2261 & w2262;
assign w2264 = pi077 & ~pi149;
assign w2265 = pi076 & ~pi148;
assign w2266 = ~w2264 & ~w2265;
assign w2267 = ~w2263 & w2266;
assign w2268 = ~pi074 & pi146;
assign w2269 = ~pi073 & pi145;
assign w2270 = ~w2268 & ~w2269;
assign w2271 = ~pi076 & pi148;
assign w2272 = ~pi075 & pi147;
assign w2273 = ~w2271 & ~w2272;
assign w2274 = w2270 & w2273;
assign w2275 = ~w2267 & w2274;
assign w2276 = pi075 & ~pi147;
assign w2277 = pi074 & ~pi146;
assign w2278 = ~w2276 & ~w2277;
assign w2279 = w2270 & ~w2278;
assign w2280 = pi073 & ~pi145;
assign w2281 = pi071 & ~pi143;
assign w2282 = pi072 & ~pi144;
assign w2283 = ~w2280 & ~w2281;
assign w2284 = ~w2282 & w2283;
assign w2285 = ~w2279 & w2284;
assign w2286 = ~w2275 & w2285;
assign w2287 = ~pi071 & pi143;
assign w2288 = ~pi072 & pi144;
assign w2289 = ~w2281 & w2288;
assign w2290 = ~w2287 & ~w2289;
assign w2291 = ~w2286 & w2290;
assign w2292 = pi078 & ~pi198;
assign w2293 = pi077 & ~pi197;
assign w2294 = ~w2292 & ~w2293;
assign w2295 = ~pi076 & pi196;
assign w2296 = ~pi077 & pi197;
assign w2297 = ~w2295 & ~w2296;
assign w2298 = ~w2294 & w2297;
assign w2299 = pi074 & ~pi194;
assign w2300 = pi073 & ~pi193;
assign w2301 = ~w2299 & ~w2300;
assign w2302 = pi076 & ~pi196;
assign w2303 = pi075 & ~pi195;
assign w2304 = ~w2302 & ~w2303;
assign w2305 = w2301 & w2304;
assign w2306 = ~w2298 & w2305;
assign w2307 = ~pi075 & pi195;
assign w2308 = ~pi074 & pi194;
assign w2309 = ~w2307 & ~w2308;
assign w2310 = w2301 & ~w2309;
assign w2311 = ~pi071 & pi191;
assign w2312 = ~pi073 & pi193;
assign w2313 = ~pi072 & pi192;
assign w2314 = ~w2311 & ~w2312;
assign w2315 = ~w2313 & w2314;
assign w2316 = ~w2310 & w2315;
assign w2317 = ~w2306 & w2316;
assign w2318 = pi071 & ~pi191;
assign w2319 = pi072 & ~pi192;
assign w2320 = ~w2311 & w2319;
assign w2321 = ~w2318 & ~w2320;
assign w2322 = ~w2317 & w2321;
assign w2323 = ~w2291 & w2322;
assign w2324 = ~w2260 & w2323;
assign w2325 = w2230 & w2324;
assign w2326 = pi078 & ~pi102;
assign w2327 = pi077 & ~pi101;
assign w2328 = ~w2326 & ~w2327;
assign w2329 = ~pi077 & pi101;
assign w2330 = ~pi076 & pi100;
assign w2331 = ~w2329 & ~w2330;
assign w2332 = ~w2328 & w2331;
assign w2333 = pi076 & ~pi100;
assign w2334 = pi075 & ~pi099;
assign w2335 = ~w2333 & ~w2334;
assign w2336 = ~pi075 & pi099;
assign w2337 = ~pi074 & pi098;
assign w2338 = ~w2336 & ~w2337;
assign w2339 = (w2338 & w2332) | (w2338 & w16211) | (w2332 & w16211);
assign w2340 = pi074 & ~pi098;
assign w2341 = pi073 & ~pi097;
assign w2342 = ~w2340 & ~w2341;
assign w2343 = ~w2339 & w2342;
assign w2344 = ~pi071 & pi095;
assign w2345 = ~pi073 & pi097;
assign w2346 = ~pi072 & pi096;
assign w2347 = ~w2345 & ~w2346;
assign w2348 = ~w2344 & w2347;
assign w2349 = ~w2343 & w2348;
assign w2350 = pi072 & ~pi096;
assign w2351 = pi071 & ~pi095;
assign w2352 = ~w2350 & ~w2351;
assign w2353 = ~w2344 & ~w2352;
assign w2354 = ~w2349 & ~w2353;
assign w2355 = ~pi077 & pi093;
assign w2356 = pi078 & ~pi094;
assign w2357 = ~w2355 & w2356;
assign w2358 = pi077 & ~pi093;
assign w2359 = pi076 & ~pi092;
assign w2360 = ~w2358 & ~w2359;
assign w2361 = ~w2357 & w2360;
assign w2362 = ~pi076 & pi092;
assign w2363 = ~pi075 & pi091;
assign w2364 = ~w2362 & ~w2363;
assign w2365 = pi075 & ~pi091;
assign w2366 = pi074 & ~pi090;
assign w2367 = ~w2365 & ~w2366;
assign w2368 = (w2367 & w2361) | (w2367 & w16212) | (w2361 & w16212);
assign w2369 = ~pi074 & pi090;
assign w2370 = ~pi073 & pi089;
assign w2371 = ~w2369 & ~w2370;
assign w2372 = ~w2368 & w2371;
assign w2373 = pi071 & ~pi087;
assign w2374 = pi072 & ~pi088;
assign w2375 = pi073 & ~pi089;
assign w2376 = ~w2373 & ~w2374;
assign w2377 = ~w2375 & w2376;
assign w2378 = ~w2372 & w2377;
assign w2379 = ~pi071 & pi087;
assign w2380 = ~pi072 & pi088;
assign w2381 = ~w2373 & w2380;
assign w2382 = ~w2379 & ~w2381;
assign w2383 = ~w2378 & w2382;
assign w2384 = w2354 & ~w2383;
assign w2385 = w2325 & w2384;
assign w2386 = w2167 & w2385;
assign w2387 = w1950 & w2386;
assign w2388 = pi075 & ~pi179;
assign w2389 = ~pi077 & pi181;
assign w2390 = pi078 & ~pi182;
assign w2391 = ~w2389 & w2390;
assign w2392 = pi077 & ~pi181;
assign w2393 = pi076 & ~pi180;
assign w2394 = ~w2392 & ~w2393;
assign w2395 = ~w2391 & w2394;
assign w2396 = ~pi076 & pi180;
assign w2397 = ~pi075 & pi179;
assign w2398 = ~w2396 & ~w2397;
assign w2399 = (~w2388 & w2395) | (~w2388 & w16213) | (w2395 & w16213);
assign w2400 = ~pi074 & pi178;
assign w2401 = ~w2399 & ~w2400;
assign w2402 = pi074 & ~pi178;
assign w2403 = pi073 & ~pi177;
assign w2404 = ~w2402 & ~w2403;
assign w2405 = ~w2401 & w2404;
assign w2406 = ~pi071 & pi175;
assign w2407 = ~pi072 & pi176;
assign w2408 = ~pi073 & pi177;
assign w2409 = ~w2406 & ~w2407;
assign w2410 = ~w2408 & w2409;
assign w2411 = ~w2405 & w2410;
assign w2412 = pi071 & ~pi175;
assign w2413 = pi072 & ~pi176;
assign w2414 = ~w2406 & w2413;
assign w2415 = ~w2412 & ~w2414;
assign w2416 = ~w2411 & w2415;
assign w2417 = ~pi071 & pi159;
assign w2418 = pi078 & ~pi166;
assign w2419 = pi077 & ~pi165;
assign w2420 = ~w2418 & ~w2419;
assign w2421 = ~pi076 & pi164;
assign w2422 = ~pi077 & pi165;
assign w2423 = ~w2421 & ~w2422;
assign w2424 = ~w2420 & w2423;
assign w2425 = pi076 & ~pi164;
assign w2426 = pi075 & ~pi163;
assign w2427 = ~w2425 & ~w2426;
assign w2428 = ~pi075 & pi163;
assign w2429 = ~pi074 & pi162;
assign w2430 = ~w2428 & ~w2429;
assign w2431 = (w2430 & w2424) | (w2430 & w16214) | (w2424 & w16214);
assign w2432 = pi074 & ~pi162;
assign w2433 = pi073 & ~pi161;
assign w2434 = ~w2432 & ~w2433;
assign w2435 = ~w2431 & w2434;
assign w2436 = ~pi072 & pi160;
assign w2437 = ~pi073 & pi161;
assign w2438 = ~w2436 & ~w2437;
assign w2439 = ~w2435 & w2438;
assign w2440 = pi071 & ~pi159;
assign w2441 = pi072 & ~pi160;
assign w2442 = ~w2440 & ~w2441;
assign w2443 = ~w2439 & w2442;
assign w2444 = ~w2417 & ~w2443;
assign w2445 = w2416 & ~w2444;
assign w2446 = pi078 & ~pi126;
assign w2447 = pi077 & ~pi125;
assign w2448 = ~w2446 & ~w2447;
assign w2449 = ~pi077 & pi125;
assign w2450 = ~pi076 & pi124;
assign w2451 = ~w2449 & ~w2450;
assign w2452 = ~w2448 & w2451;
assign w2453 = pi076 & ~pi124;
assign w2454 = pi075 & ~pi123;
assign w2455 = ~w2453 & ~w2454;
assign w2456 = ~pi075 & pi123;
assign w2457 = ~pi074 & pi122;
assign w2458 = ~w2456 & ~w2457;
assign w2459 = (w2458 & w2452) | (w2458 & w16215) | (w2452 & w16215);
assign w2460 = pi074 & ~pi122;
assign w2461 = pi073 & ~pi121;
assign w2462 = ~w2460 & ~w2461;
assign w2463 = ~w2459 & w2462;
assign w2464 = ~pi073 & pi121;
assign w2465 = ~pi072 & pi120;
assign w2466 = ~w2464 & ~w2465;
assign w2467 = ~w2463 & w2466;
assign w2468 = pi072 & ~pi120;
assign w2469 = pi071 & ~pi119;
assign w2470 = ~w2468 & ~w2469;
assign w2471 = ~w2467 & w2470;
assign w2472 = ~pi071 & pi119;
assign w2473 = ~w2471 & ~w2472;
assign w2474 = ~pi071 & pi103;
assign w2475 = pi073 & ~pi105;
assign w2476 = pi078 & ~pi110;
assign w2477 = pi077 & ~pi109;
assign w2478 = ~w2476 & ~w2477;
assign w2479 = ~pi077 & pi109;
assign w2480 = ~pi076 & pi108;
assign w2481 = ~w2479 & ~w2480;
assign w2482 = ~w2478 & w2481;
assign w2483 = pi074 & ~pi106;
assign w2484 = pi076 & ~pi108;
assign w2485 = pi075 & ~pi107;
assign w2486 = ~w2483 & ~w2484;
assign w2487 = ~w2485 & w2486;
assign w2488 = ~w2482 & w2487;
assign w2489 = ~pi073 & pi105;
assign w2490 = ~pi074 & pi106;
assign w2491 = ~pi075 & pi107;
assign w2492 = ~w2483 & w2491;
assign w2493 = ~w2489 & ~w2490;
assign w2494 = ~w2492 & w2493;
assign w2495 = (~w2475 & w2488) | (~w2475 & w16216) | (w2488 & w16216);
assign w2496 = ~pi072 & pi104;
assign w2497 = ~w2495 & ~w2496;
assign w2498 = pi072 & ~pi104;
assign w2499 = pi071 & ~pi103;
assign w2500 = ~w2498 & ~w2499;
assign w2501 = ~w2497 & w2500;
assign w2502 = ~w2474 & ~w2501;
assign w2503 = ~w2473 & ~w2502;
assign w2504 = w2445 & w2503;
assign w2505 = pi075 & ~pi083;
assign w2506 = pi076 & ~pi084;
assign w2507 = ~pi076 & pi084;
assign w2508 = pi077 & ~pi085;
assign w2509 = pi078 & ~pi086;
assign w2510 = ~w2508 & ~w2509;
assign w2511 = ~pi077 & pi085;
assign w2512 = ~w2507 & ~w2511;
assign w2513 = ~w2510 & w2512;
assign w2514 = ~w2505 & ~w2506;
assign w2515 = ~w2513 & w2514;
assign w2516 = ~pi074 & pi082;
assign w2517 = ~pi073 & pi081;
assign w2518 = ~pi072 & pi080;
assign w2519 = ~w2517 & ~w2518;
assign w2520 = ~pi075 & pi083;
assign w2521 = ~w2516 & ~w2520;
assign w2522 = w2519 & w2521;
assign w2523 = ~w2515 & w2522;
assign w2524 = pi071 & ~pi079;
assign w2525 = pi074 & ~pi082;
assign w2526 = pi073 & ~pi081;
assign w2527 = ~w2525 & ~w2526;
assign w2528 = w2519 & ~w2527;
assign w2529 = pi072 & ~pi080;
assign w2530 = ~w2524 & ~w2529;
assign w2531 = ~w2528 & w2530;
assign w2532 = ~w2523 & w2531;
assign w2533 = ~pi071 & pi079;
assign w2534 = ~w2532 & ~w2533;
assign w2535 = w955 & ~w2534;
assign w2536 = w2504 & w2535;
assign w2537 = w2387 & w2536;
assign w2538 = ~w1767 & w2537;
assign w2539 = (~w1230 & ~w1423) | (~w1230 & w16217) | (~w1423 & w16217);
assign w2540 = w2538 & ~w2539;
assign w2541 = pi005 & w2540;
assign w2542 = ~w950 & ~w1198;
assign w2543 = ~w2532 & w2542;
assign w2544 = ~w367 & w16218;
assign w2545 = w347 & ~w2544;
assign w2546 = w922 & ~w2545;
assign w2547 = w2543 & w2546;
assign w2548 = ~w344 & w952;
assign w2549 = ~w951 & ~w1170;
assign w2550 = ~w2533 & w2549;
assign w2551 = w2548 & w2550;
assign w2552 = w2547 & w2551;
assign w2553 = pi006 & w2552;
assign w2554 = w29 & w467;
assign w2555 = ~w918 & ~w2554;
assign w2556 = w1670 & w1756;
assign w2557 = ~w955 & w1420;
assign w2558 = w1419 & ~w2557;
assign w2559 = w1298 & w2558;
assign w2560 = w2556 & w2559;
assign w2561 = ~w2555 & w2560;
assign w2562 = ~w1759 & w2561;
assign w2563 = pi003 & w2562;
assign w2564 = (w467 & ~w1423) | (w467 & w16219) | (~w1423 & w16219);
assign w2565 = w437 & ~w955;
assign w2566 = w406 & ~w2565;
assign w2567 = w280 & w2566;
assign w2568 = w917 & w2567;
assign w2569 = ~w469 & w2568;
assign w2570 = ~w2564 & w2569;
assign w2571 = pi001 & w2570;
assign w2572 = w437 & w1421;
assign w2573 = ~w918 & ~w2572;
assign w2574 = (~w1420 & ~w1423) | (~w1420 & w16220) | (~w1423 & w16220);
assign w2575 = ~w2573 & ~w2574;
assign w2576 = pi004 & w2575;
assign w2577 = ~w2541 & ~w2553;
assign w2578 = ~w2563 & ~w2571;
assign w2579 = ~w2576 & w2578;
assign w2580 = w2577 & w2579;
assign w2581 = ~w918 & w16221;
assign w2582 = ~w2574 & ~w2581;
assign w2583 = w373 & ~w918;
assign w2584 = ~w2570 & w2583;
assign w2585 = w2582 & ~w2584;
assign w2586 = (~w2534 & ~w2538) | (~w2534 & w16222) | (~w2538 & w16222);
assign w2587 = ~w1199 & ~w2561;
assign w2588 = ~w2586 & ~w2587;
assign w2589 = w2585 & w2588;
assign w2590 = ~w2552 & w2589;
assign w2591 = pi006 & w2590;
assign w2592 = ~pi087 & pi095;
assign w2593 = ~w2344 & ~w2533;
assign w2594 = ~w2592 & w2593;
assign w2595 = ~w281 & ~w957;
assign w2596 = w2594 & w2595;
assign w2597 = w2551 & w2596;
assign w2598 = pi091 & ~pi099;
assign w2599 = pi092 & ~pi100;
assign w2600 = ~pi092 & pi100;
assign w2601 = pi094 & ~pi102;
assign w2602 = pi093 & ~pi101;
assign w2603 = ~w2601 & ~w2602;
assign w2604 = ~pi093 & pi101;
assign w2605 = ~w2600 & ~w2604;
assign w2606 = ~w2603 & w2605;
assign w2607 = ~w2598 & ~w2599;
assign w2608 = ~w2606 & w2607;
assign w2609 = ~pi091 & pi099;
assign w2610 = ~pi090 & pi098;
assign w2611 = ~w2609 & ~w2610;
assign w2612 = ~w2608 & w2611;
assign w2613 = pi090 & ~pi098;
assign w2614 = pi089 & ~pi097;
assign w2615 = ~w2613 & ~w2614;
assign w2616 = ~w2612 & w2615;
assign w2617 = ~pi089 & pi097;
assign w2618 = ~pi088 & pi096;
assign w2619 = ~w2617 & ~w2618;
assign w2620 = ~w2616 & w2619;
assign w2621 = pi088 & ~pi096;
assign w2622 = pi087 & ~pi095;
assign w2623 = ~w2621 & ~w2622;
assign w2624 = ~w2620 & w2623;
assign w2625 = ~w2343 & w2347;
assign w2626 = w2352 & ~w2625;
assign w2627 = ~w2624 & ~w2626;
assign w2628 = w2543 & w2627;
assign w2629 = w310 & w2546;
assign w2630 = w2597 & w2629;
assign w2631 = w2628 & w2630;
assign w2632 = ~w983 & w2631;
assign w2633 = pi008 & w2632;
assign w2634 = ~w918 & ~w2570;
assign w2635 = w2561 & ~w2634;
assign w2636 = pi004 & w2635;
assign w2637 = (~w2383 & ~w2538) | (~w2383 & w16223) | (~w2538 & w16223);
assign w2638 = w1012 & ~w2561;
assign w2639 = pi087 & ~pi103;
assign w2640 = pi089 & ~pi105;
assign w2641 = pi088 & ~pi104;
assign w2642 = ~pi089 & pi105;
assign w2643 = ~pi090 & pi106;
assign w2644 = pi091 & ~pi107;
assign w2645 = pi090 & ~pi106;
assign w2646 = pi092 & ~pi108;
assign w2647 = pi093 & ~pi109;
assign w2648 = ~pi093 & pi109;
assign w2649 = pi094 & ~pi110;
assign w2650 = ~w2648 & w2649;
assign w2651 = ~w2646 & ~w2647;
assign w2652 = ~w2650 & w2651;
assign w2653 = ~pi092 & pi108;
assign w2654 = ~pi091 & pi107;
assign w2655 = ~w2653 & ~w2654;
assign w2656 = ~w2652 & w2655;
assign w2657 = ~w2644 & ~w2645;
assign w2658 = ~w2656 & w2657;
assign w2659 = ~w2642 & ~w2643;
assign w2660 = ~w2658 & w2659;
assign w2661 = ~w2640 & ~w2641;
assign w2662 = ~w2660 & w2661;
assign w2663 = ~pi088 & pi104;
assign w2664 = ~pi087 & pi103;
assign w2665 = ~w2663 & ~w2664;
assign w2666 = ~w2662 & w2665;
assign w2667 = ~w2639 & ~w2666;
assign w2668 = ~pi087 & pi159;
assign w2669 = pi092 & ~pi164;
assign w2670 = pi091 & ~pi163;
assign w2671 = ~pi092 & pi164;
assign w2672 = pi093 & ~pi165;
assign w2673 = ~pi093 & pi165;
assign w2674 = pi094 & ~pi166;
assign w2675 = ~w2673 & w2674;
assign w2676 = (~w2671 & w2675) | (~w2671 & w16224) | (w2675 & w16224);
assign w2677 = ~w2669 & ~w2670;
assign w2678 = ~w2676 & w2677;
assign w2679 = ~pi090 & pi162;
assign w2680 = ~pi091 & pi163;
assign w2681 = ~w2679 & ~w2680;
assign w2682 = ~w2678 & w2681;
assign w2683 = pi090 & ~pi162;
assign w2684 = pi089 & ~pi161;
assign w2685 = ~w2683 & ~w2684;
assign w2686 = ~w2682 & w2685;
assign w2687 = ~pi089 & pi161;
assign w2688 = ~pi088 & pi160;
assign w2689 = ~w2687 & ~w2688;
assign w2690 = ~w2686 & w2689;
assign w2691 = pi087 & ~pi159;
assign w2692 = pi088 & ~pi160;
assign w2693 = ~w2691 & ~w2692;
assign w2694 = ~w2690 & w2693;
assign w2695 = ~w2668 & ~w2694;
assign w2696 = ~pi087 & pi175;
assign w2697 = pi092 & ~pi180;
assign w2698 = pi091 & ~pi179;
assign w2699 = ~pi092 & pi180;
assign w2700 = pi093 & ~pi181;
assign w2701 = ~pi093 & pi181;
assign w2702 = pi094 & ~pi182;
assign w2703 = ~w2701 & w2702;
assign w2704 = (~w2699 & w2703) | (~w2699 & w16225) | (w2703 & w16225);
assign w2705 = ~w2697 & ~w2698;
assign w2706 = ~w2704 & w2705;
assign w2707 = ~pi090 & pi178;
assign w2708 = ~pi091 & pi179;
assign w2709 = ~w2707 & ~w2708;
assign w2710 = ~w2706 & w2709;
assign w2711 = pi090 & ~pi178;
assign w2712 = pi089 & ~pi177;
assign w2713 = ~w2711 & ~w2712;
assign w2714 = ~w2710 & w2713;
assign w2715 = ~pi089 & pi177;
assign w2716 = ~pi088 & pi176;
assign w2717 = ~w2715 & ~w2716;
assign w2718 = ~w2714 & w2717;
assign w2719 = pi087 & ~pi175;
assign w2720 = pi088 & ~pi176;
assign w2721 = ~w2719 & ~w2720;
assign w2722 = ~w2718 & w2721;
assign w2723 = ~w2696 & ~w2722;
assign w2724 = ~w2695 & ~w2723;
assign w2725 = pi087 & ~pi119;
assign w2726 = ~pi087 & pi119;
assign w2727 = ~pi088 & pi120;
assign w2728 = pi088 & ~pi120;
assign w2729 = pi089 & ~pi121;
assign w2730 = ~pi090 & pi122;
assign w2731 = ~pi089 & pi121;
assign w2732 = pi091 & ~pi123;
assign w2733 = pi090 & ~pi122;
assign w2734 = ~pi092 & pi124;
assign w2735 = ~pi091 & pi123;
assign w2736 = pi092 & ~pi124;
assign w2737 = pi093 & ~pi125;
assign w2738 = ~pi093 & pi125;
assign w2739 = pi094 & ~pi126;
assign w2740 = ~w2738 & w2739;
assign w2741 = ~w2736 & ~w2737;
assign w2742 = ~w2740 & w2741;
assign w2743 = ~w2734 & ~w2735;
assign w2744 = ~w2742 & w2743;
assign w2745 = ~w2732 & ~w2733;
assign w2746 = ~w2744 & w2745;
assign w2747 = ~w2730 & ~w2731;
assign w2748 = ~w2746 & w2747;
assign w2749 = ~w2728 & ~w2729;
assign w2750 = ~w2748 & w2749;
assign w2751 = ~w2726 & ~w2727;
assign w2752 = ~w2750 & w2751;
assign w2753 = ~w2725 & ~w2752;
assign w2754 = w2724 & w2753;
assign w2755 = w2667 & w2754;
assign w2756 = ~pi087 & pi223;
assign w2757 = ~pi089 & pi225;
assign w2758 = ~pi088 & pi224;
assign w2759 = pi089 & ~pi225;
assign w2760 = pi090 & ~pi226;
assign w2761 = ~pi090 & pi226;
assign w2762 = ~pi091 & pi227;
assign w2763 = pi092 & ~pi228;
assign w2764 = pi091 & ~pi227;
assign w2765 = pi093 & ~pi229;
assign w2766 = pi094 & ~pi230;
assign w2767 = ~w2765 & ~w2766;
assign w2768 = ~pi092 & pi228;
assign w2769 = ~pi093 & pi229;
assign w2770 = ~w2768 & ~w2769;
assign w2771 = ~w2767 & w2770;
assign w2772 = ~w2763 & ~w2764;
assign w2773 = ~w2771 & w2772;
assign w2774 = ~w2761 & ~w2762;
assign w2775 = ~w2773 & w2774;
assign w2776 = ~w2759 & ~w2760;
assign w2777 = ~w2775 & w2776;
assign w2778 = ~w2757 & ~w2758;
assign w2779 = ~w2777 & w2778;
assign w2780 = pi088 & ~pi224;
assign w2781 = pi087 & ~pi223;
assign w2782 = ~w2780 & ~w2781;
assign w2783 = ~w2779 & w2782;
assign w2784 = ~w2756 & ~w2783;
assign w2785 = ~pi087 & pi263;
assign w2786 = pi092 & ~pi268;
assign w2787 = pi091 & ~pi267;
assign w2788 = ~pi092 & pi268;
assign w2789 = pi093 & ~pi269;
assign w2790 = pi094 & ~pi270;
assign w2791 = ~w2789 & ~w2790;
assign w2792 = ~pi093 & pi269;
assign w2793 = ~w2788 & ~w2792;
assign w2794 = ~w2791 & w2793;
assign w2795 = ~w2786 & ~w2787;
assign w2796 = ~w2794 & w2795;
assign w2797 = ~pi091 & pi267;
assign w2798 = ~pi090 & pi266;
assign w2799 = ~w2797 & ~w2798;
assign w2800 = ~w2796 & w2799;
assign w2801 = pi090 & ~pi266;
assign w2802 = pi089 & ~pi265;
assign w2803 = ~w2801 & ~w2802;
assign w2804 = ~w2800 & w2803;
assign w2805 = ~pi089 & pi265;
assign w2806 = ~pi088 & pi264;
assign w2807 = ~w2805 & ~w2806;
assign w2808 = ~w2804 & w2807;
assign w2809 = pi088 & ~pi264;
assign w2810 = pi087 & ~pi263;
assign w2811 = ~w2809 & ~w2810;
assign w2812 = ~w2808 & w2811;
assign w2813 = ~w2785 & ~w2812;
assign w2814 = ~pi087 & pi247;
assign w2815 = pi092 & ~pi252;
assign w2816 = pi091 & ~pi251;
assign w2817 = ~pi092 & pi252;
assign w2818 = pi093 & ~pi253;
assign w2819 = pi094 & ~pi254;
assign w2820 = ~w2818 & ~w2819;
assign w2821 = ~pi093 & pi253;
assign w2822 = ~w2817 & ~w2821;
assign w2823 = ~w2820 & w2822;
assign w2824 = ~w2815 & ~w2816;
assign w2825 = ~w2823 & w2824;
assign w2826 = ~pi091 & pi251;
assign w2827 = ~pi090 & pi250;
assign w2828 = ~w2826 & ~w2827;
assign w2829 = ~w2825 & w2828;
assign w2830 = pi090 & ~pi250;
assign w2831 = pi089 & ~pi249;
assign w2832 = ~w2830 & ~w2831;
assign w2833 = ~w2829 & w2832;
assign w2834 = ~pi089 & pi249;
assign w2835 = ~pi088 & pi248;
assign w2836 = ~w2834 & ~w2835;
assign w2837 = ~w2833 & w2836;
assign w2838 = pi088 & ~pi248;
assign w2839 = pi087 & ~pi247;
assign w2840 = ~w2838 & ~w2839;
assign w2841 = ~w2837 & w2840;
assign w2842 = ~w2814 & ~w2841;
assign w2843 = ~w2813 & ~w2842;
assign w2844 = ~w2784 & w2843;
assign w2845 = ~pi087 & pi151;
assign w2846 = pi092 & ~pi156;
assign w2847 = pi091 & ~pi155;
assign w2848 = ~pi092 & pi156;
assign w2849 = pi093 & ~pi157;
assign w2850 = pi094 & ~pi158;
assign w2851 = ~w2849 & ~w2850;
assign w2852 = ~pi093 & pi157;
assign w2853 = ~w2848 & ~w2852;
assign w2854 = ~w2851 & w2853;
assign w2855 = ~w2846 & ~w2847;
assign w2856 = ~w2854 & w2855;
assign w2857 = ~pi091 & pi155;
assign w2858 = ~pi090 & pi154;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = ~w2856 & w2859;
assign w2861 = pi090 & ~pi154;
assign w2862 = pi089 & ~pi153;
assign w2863 = ~w2861 & ~w2862;
assign w2864 = ~w2860 & w2863;
assign w2865 = ~pi089 & pi153;
assign w2866 = ~pi088 & pi152;
assign w2867 = ~w2865 & ~w2866;
assign w2868 = ~w2864 & w2867;
assign w2869 = pi088 & ~pi152;
assign w2870 = pi087 & ~pi151;
assign w2871 = ~w2869 & ~w2870;
assign w2872 = ~w2868 & w2871;
assign w2873 = ~w2845 & ~w2872;
assign w2874 = ~pi087 & pi199;
assign w2875 = pi093 & ~pi205;
assign w2876 = pi094 & ~pi206;
assign w2877 = ~w2875 & ~w2876;
assign w2878 = ~pi093 & pi205;
assign w2879 = ~pi092 & pi204;
assign w2880 = ~w2878 & ~w2879;
assign w2881 = ~w2877 & w2880;
assign w2882 = pi091 & ~pi203;
assign w2883 = pi092 & ~pi204;
assign w2884 = ~w2882 & ~w2883;
assign w2885 = ~w2881 & w2884;
assign w2886 = ~pi091 & pi203;
assign w2887 = ~pi090 & pi202;
assign w2888 = ~w2886 & ~w2887;
assign w2889 = ~w2885 & w2888;
assign w2890 = pi090 & ~pi202;
assign w2891 = pi089 & ~pi201;
assign w2892 = ~w2890 & ~w2891;
assign w2893 = ~w2889 & w2892;
assign w2894 = ~pi089 & pi201;
assign w2895 = ~pi088 & pi200;
assign w2896 = ~w2894 & ~w2895;
assign w2897 = ~w2893 & w2896;
assign w2898 = pi088 & ~pi200;
assign w2899 = pi087 & ~pi199;
assign w2900 = ~w2898 & ~w2899;
assign w2901 = ~w2897 & w2900;
assign w2902 = ~w2874 & ~w2901;
assign w2903 = ~pi087 & pi207;
assign w2904 = pi093 & ~pi213;
assign w2905 = pi094 & ~pi214;
assign w2906 = ~w2904 & ~w2905;
assign w2907 = ~pi093 & pi213;
assign w2908 = ~pi092 & pi212;
assign w2909 = ~w2907 & ~w2908;
assign w2910 = ~w2906 & w2909;
assign w2911 = pi091 & ~pi211;
assign w2912 = pi092 & ~pi212;
assign w2913 = ~w2911 & ~w2912;
assign w2914 = ~w2910 & w2913;
assign w2915 = ~pi091 & pi211;
assign w2916 = ~pi090 & pi210;
assign w2917 = ~w2915 & ~w2916;
assign w2918 = ~w2914 & w2917;
assign w2919 = pi090 & ~pi210;
assign w2920 = pi089 & ~pi209;
assign w2921 = ~w2919 & ~w2920;
assign w2922 = ~w2918 & w2921;
assign w2923 = ~pi089 & pi209;
assign w2924 = ~pi088 & pi208;
assign w2925 = ~w2923 & ~w2924;
assign w2926 = ~w2922 & w2925;
assign w2927 = pi088 & ~pi208;
assign w2928 = pi087 & ~pi207;
assign w2929 = ~w2927 & ~w2928;
assign w2930 = ~w2926 & w2929;
assign w2931 = ~w2903 & ~w2930;
assign w2932 = ~w2902 & ~w2931;
assign w2933 = ~pi087 & pi167;
assign w2934 = pi093 & ~pi173;
assign w2935 = pi094 & ~pi174;
assign w2936 = ~w2934 & ~w2935;
assign w2937 = ~pi092 & pi172;
assign w2938 = ~pi093 & pi173;
assign w2939 = ~w2937 & ~w2938;
assign w2940 = ~w2936 & w2939;
assign w2941 = pi091 & ~pi171;
assign w2942 = pi092 & ~pi172;
assign w2943 = ~w2941 & ~w2942;
assign w2944 = ~w2940 & w2943;
assign w2945 = ~pi090 & pi170;
assign w2946 = ~pi091 & pi171;
assign w2947 = ~w2945 & ~w2946;
assign w2948 = ~w2944 & w2947;
assign w2949 = pi090 & ~pi170;
assign w2950 = pi089 & ~pi169;
assign w2951 = ~w2949 & ~w2950;
assign w2952 = ~w2948 & w2951;
assign w2953 = ~pi089 & pi169;
assign w2954 = ~pi088 & pi168;
assign w2955 = ~w2953 & ~w2954;
assign w2956 = ~w2952 & w2955;
assign w2957 = pi088 & ~pi168;
assign w2958 = pi087 & ~pi167;
assign w2959 = ~w2957 & ~w2958;
assign w2960 = ~w2956 & w2959;
assign w2961 = ~w2933 & ~w2960;
assign w2962 = pi093 & ~pi133;
assign w2963 = pi094 & ~pi134;
assign w2964 = ~w2962 & ~w2963;
assign w2965 = ~pi093 & pi133;
assign w2966 = ~pi092 & pi132;
assign w2967 = ~w2965 & ~w2966;
assign w2968 = ~w2964 & w2967;
assign w2969 = pi092 & ~pi132;
assign w2970 = pi091 & ~pi131;
assign w2971 = ~w2969 & ~w2970;
assign w2972 = ~w2968 & w2971;
assign w2973 = ~pi091 & pi131;
assign w2974 = ~pi090 & pi130;
assign w2975 = ~w2973 & ~w2974;
assign w2976 = ~w2972 & w2975;
assign w2977 = pi090 & ~pi130;
assign w2978 = pi089 & ~pi129;
assign w2979 = ~w2977 & ~w2978;
assign w2980 = ~w2976 & w2979;
assign w2981 = ~pi089 & pi129;
assign w2982 = ~pi088 & pi128;
assign w2983 = ~w2981 & ~w2982;
assign w2984 = ~w2980 & w2983;
assign w2985 = pi088 & ~pi128;
assign w2986 = pi087 & ~pi127;
assign w2987 = ~w2985 & ~w2986;
assign w2988 = ~w2984 & w2987;
assign w2989 = ~pi087 & pi127;
assign w2990 = ~w2988 & ~w2989;
assign w2991 = pi087 & ~pi191;
assign w2992 = ~pi093 & pi197;
assign w2993 = pi094 & ~pi198;
assign w2994 = ~w2992 & w2993;
assign w2995 = pi093 & ~pi197;
assign w2996 = pi092 & ~pi196;
assign w2997 = ~w2995 & ~w2996;
assign w2998 = ~w2994 & w2997;
assign w2999 = ~pi092 & pi196;
assign w3000 = ~pi091 & pi195;
assign w3001 = ~w2999 & ~w3000;
assign w3002 = ~w2998 & w3001;
assign w3003 = pi091 & ~pi195;
assign w3004 = pi090 & ~pi194;
assign w3005 = ~w3003 & ~w3004;
assign w3006 = ~w3002 & w3005;
assign w3007 = ~pi090 & pi194;
assign w3008 = ~pi089 & pi193;
assign w3009 = ~w3007 & ~w3008;
assign w3010 = ~w3006 & w3009;
assign w3011 = pi089 & ~pi193;
assign w3012 = pi088 & ~pi192;
assign w3013 = ~w3011 & ~w3012;
assign w3014 = ~w3010 & w3013;
assign w3015 = ~pi087 & pi191;
assign w3016 = ~pi088 & pi192;
assign w3017 = ~w3015 & ~w3016;
assign w3018 = ~w3014 & w3017;
assign w3019 = ~w2991 & ~w3018;
assign w3020 = pi087 & ~pi143;
assign w3021 = ~pi093 & pi149;
assign w3022 = pi094 & ~pi150;
assign w3023 = ~w3021 & w3022;
assign w3024 = pi093 & ~pi149;
assign w3025 = pi092 & ~pi148;
assign w3026 = ~w3024 & ~w3025;
assign w3027 = ~w3023 & w3026;
assign w3028 = ~pi092 & pi148;
assign w3029 = ~pi091 & pi147;
assign w3030 = ~w3028 & ~w3029;
assign w3031 = ~w3027 & w3030;
assign w3032 = pi091 & ~pi147;
assign w3033 = pi090 & ~pi146;
assign w3034 = ~w3032 & ~w3033;
assign w3035 = ~w3031 & w3034;
assign w3036 = ~pi090 & pi146;
assign w3037 = ~pi089 & pi145;
assign w3038 = ~w3036 & ~w3037;
assign w3039 = ~w3035 & w3038;
assign w3040 = pi089 & ~pi145;
assign w3041 = pi088 & ~pi144;
assign w3042 = ~w3040 & ~w3041;
assign w3043 = ~w3039 & w3042;
assign w3044 = ~pi087 & pi143;
assign w3045 = ~pi088 & pi144;
assign w3046 = ~w3044 & ~w3045;
assign w3047 = ~w3043 & w3046;
assign w3048 = ~w3020 & ~w3047;
assign w3049 = w3019 & w3048;
assign w3050 = ~w2873 & ~w2961;
assign w3051 = ~w2990 & w3050;
assign w3052 = w2932 & w3049;
assign w3053 = w3051 & w3052;
assign w3054 = w2844 & w3053;
assign w3055 = ~pi087 & pi239;
assign w3056 = pi094 & ~pi246;
assign w3057 = pi093 & ~pi245;
assign w3058 = ~w3056 & ~w3057;
assign w3059 = ~pi093 & pi245;
assign w3060 = ~pi092 & pi244;
assign w3061 = ~w3059 & ~w3060;
assign w3062 = ~w3058 & w3061;
assign w3063 = pi092 & ~pi244;
assign w3064 = pi091 & ~pi243;
assign w3065 = ~w3063 & ~w3064;
assign w3066 = ~pi091 & pi243;
assign w3067 = ~pi090 & pi242;
assign w3068 = ~w3066 & ~w3067;
assign w3069 = (w3068 & w3062) | (w3068 & w16226) | (w3062 & w16226);
assign w3070 = pi090 & ~pi242;
assign w3071 = pi089 & ~pi241;
assign w3072 = ~w3070 & ~w3071;
assign w3073 = ~w3069 & w3072;
assign w3074 = ~pi089 & pi241;
assign w3075 = ~pi088 & pi240;
assign w3076 = ~w3074 & ~w3075;
assign w3077 = ~w3073 & w3076;
assign w3078 = pi088 & ~pi240;
assign w3079 = pi087 & ~pi239;
assign w3080 = ~w3078 & ~w3079;
assign w3081 = ~w3077 & w3080;
assign w3082 = ~w3055 & ~w3081;
assign w3083 = pi094 & ~pi238;
assign w3084 = pi093 & ~pi237;
assign w3085 = ~w3083 & ~w3084;
assign w3086 = ~pi093 & pi237;
assign w3087 = ~pi092 & pi236;
assign w3088 = ~w3086 & ~w3087;
assign w3089 = ~w3085 & w3088;
assign w3090 = pi092 & ~pi236;
assign w3091 = pi091 & ~pi235;
assign w3092 = ~w3090 & ~w3091;
assign w3093 = ~pi091 & pi235;
assign w3094 = ~pi090 & pi234;
assign w3095 = ~w3093 & ~w3094;
assign w3096 = (w3095 & w3089) | (w3095 & w16227) | (w3089 & w16227);
assign w3097 = pi090 & ~pi234;
assign w3098 = pi089 & ~pi233;
assign w3099 = ~w3097 & ~w3098;
assign w3100 = ~w3096 & w3099;
assign w3101 = ~pi089 & pi233;
assign w3102 = ~pi088 & pi232;
assign w3103 = ~w3101 & ~w3102;
assign w3104 = ~w3100 & w3103;
assign w3105 = pi088 & ~pi232;
assign w3106 = pi087 & ~pi231;
assign w3107 = ~w3105 & ~w3106;
assign w3108 = ~w3104 & w3107;
assign w3109 = ~pi087 & pi231;
assign w3110 = ~w3108 & ~w3109;
assign w3111 = ~w3082 & ~w3110;
assign w3112 = pi094 & ~pi262;
assign w3113 = pi093 & ~pi261;
assign w3114 = ~w3112 & ~w3113;
assign w3115 = ~pi093 & pi261;
assign w3116 = ~pi092 & pi260;
assign w3117 = ~w3115 & ~w3116;
assign w3118 = ~w3114 & w3117;
assign w3119 = pi092 & ~pi260;
assign w3120 = pi091 & ~pi259;
assign w3121 = ~w3119 & ~w3120;
assign w3122 = ~pi091 & pi259;
assign w3123 = ~pi090 & pi258;
assign w3124 = ~w3122 & ~w3123;
assign w3125 = (w3124 & w3118) | (w3124 & w16228) | (w3118 & w16228);
assign w3126 = pi090 & ~pi258;
assign w3127 = pi089 & ~pi257;
assign w3128 = ~w3126 & ~w3127;
assign w3129 = ~w3125 & w3128;
assign w3130 = ~pi089 & pi257;
assign w3131 = ~pi088 & pi256;
assign w3132 = ~w3130 & ~w3131;
assign w3133 = ~w3129 & w3132;
assign w3134 = pi088 & ~pi256;
assign w3135 = pi087 & ~pi255;
assign w3136 = ~w3134 & ~w3135;
assign w3137 = ~w3133 & w3136;
assign w3138 = ~pi087 & pi255;
assign w3139 = ~w3137 & ~w3138;
assign w3140 = pi094 & ~pi222;
assign w3141 = pi093 & ~pi221;
assign w3142 = ~w3140 & ~w3141;
assign w3143 = ~pi093 & pi221;
assign w3144 = ~pi092 & pi220;
assign w3145 = ~w3143 & ~w3144;
assign w3146 = ~w3142 & w3145;
assign w3147 = pi092 & ~pi220;
assign w3148 = pi091 & ~pi219;
assign w3149 = ~w3147 & ~w3148;
assign w3150 = ~pi091 & pi219;
assign w3151 = ~pi090 & pi218;
assign w3152 = ~w3150 & ~w3151;
assign w3153 = (w3152 & w3146) | (w3152 & w16229) | (w3146 & w16229);
assign w3154 = pi090 & ~pi218;
assign w3155 = pi089 & ~pi217;
assign w3156 = ~w3154 & ~w3155;
assign w3157 = ~w3153 & w3156;
assign w3158 = ~pi089 & pi217;
assign w3159 = ~pi088 & pi216;
assign w3160 = ~w3158 & ~w3159;
assign w3161 = ~w3157 & w3160;
assign w3162 = pi088 & ~pi216;
assign w3163 = pi087 & ~pi215;
assign w3164 = ~w3162 & ~w3163;
assign w3165 = ~w3161 & w3164;
assign w3166 = ~pi087 & pi215;
assign w3167 = ~w3165 & ~w3166;
assign w3168 = ~w3139 & ~w3167;
assign w3169 = w3111 & w3168;
assign w3170 = pi092 & ~pi140;
assign w3171 = pi091 & ~pi139;
assign w3172 = ~pi093 & pi141;
assign w3173 = pi094 & ~pi142;
assign w3174 = pi093 & ~pi141;
assign w3175 = ~w3173 & ~w3174;
assign w3176 = ~pi092 & pi140;
assign w3177 = ~w3172 & ~w3176;
assign w3178 = ~w3175 & w3177;
assign w3179 = ~w3170 & ~w3171;
assign w3180 = ~pi091 & pi139;
assign w3181 = ~pi090 & pi138;
assign w3182 = ~w3180 & ~w3181;
assign w3183 = (w3182 & w3178) | (w3182 & w16230) | (w3178 & w16230);
assign w3184 = pi090 & ~pi138;
assign w3185 = pi089 & ~pi137;
assign w3186 = ~w3184 & ~w3185;
assign w3187 = ~w3183 & w3186;
assign w3188 = ~pi089 & pi137;
assign w3189 = ~pi088 & pi136;
assign w3190 = ~w3188 & ~w3189;
assign w3191 = ~w3187 & w3190;
assign w3192 = pi088 & ~pi136;
assign w3193 = pi087 & ~pi135;
assign w3194 = ~w3192 & ~w3193;
assign w3195 = ~w3191 & w3194;
assign w3196 = ~pi087 & pi135;
assign w3197 = ~w3195 & ~w3196;
assign w3198 = pi094 & ~pi190;
assign w3199 = pi093 & ~pi189;
assign w3200 = ~w3198 & ~w3199;
assign w3201 = ~pi093 & pi189;
assign w3202 = ~pi092 & pi188;
assign w3203 = ~w3201 & ~w3202;
assign w3204 = ~w3200 & w3203;
assign w3205 = pi092 & ~pi188;
assign w3206 = pi091 & ~pi187;
assign w3207 = ~w3205 & ~w3206;
assign w3208 = ~pi091 & pi187;
assign w3209 = ~pi090 & pi186;
assign w3210 = ~w3208 & ~w3209;
assign w3211 = (w3210 & w3204) | (w3210 & w16231) | (w3204 & w16231);
assign w3212 = pi090 & ~pi186;
assign w3213 = pi089 & ~pi185;
assign w3214 = ~w3212 & ~w3213;
assign w3215 = ~w3211 & w3214;
assign w3216 = ~pi089 & pi185;
assign w3217 = ~pi088 & pi184;
assign w3218 = ~w3216 & ~w3217;
assign w3219 = ~w3215 & w3218;
assign w3220 = pi088 & ~pi184;
assign w3221 = pi087 & ~pi183;
assign w3222 = ~w3220 & ~w3221;
assign w3223 = ~w3219 & w3222;
assign w3224 = ~pi087 & pi183;
assign w3225 = ~w3223 & ~w3224;
assign w3226 = pi094 & ~pi278;
assign w3227 = pi093 & ~pi277;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = ~pi092 & pi276;
assign w3230 = ~pi093 & pi277;
assign w3231 = ~w3229 & ~w3230;
assign w3232 = ~w3228 & w3231;
assign w3233 = pi092 & ~pi276;
assign w3234 = pi091 & ~pi275;
assign w3235 = ~w3233 & ~w3234;
assign w3236 = ~w3232 & w3235;
assign w3237 = ~pi091 & pi275;
assign w3238 = ~pi090 & pi274;
assign w3239 = ~w3237 & ~w3238;
assign w3240 = ~w3236 & w3239;
assign w3241 = pi090 & ~pi274;
assign w3242 = pi089 & ~pi273;
assign w3243 = ~w3241 & ~w3242;
assign w3244 = ~w3240 & w3243;
assign w3245 = ~pi089 & pi273;
assign w3246 = ~pi088 & pi272;
assign w3247 = ~w3245 & ~w3246;
assign w3248 = ~w3244 & w3247;
assign w3249 = pi088 & ~pi272;
assign w3250 = pi087 & ~pi271;
assign w3251 = ~w3249 & ~w3250;
assign w3252 = ~w3248 & w3251;
assign w3253 = ~pi087 & pi271;
assign w3254 = ~w3252 & ~w3253;
assign w3255 = ~w3197 & ~w3225;
assign w3256 = ~w3254 & w3255;
assign w3257 = w3169 & w3256;
assign w3258 = ~w2592 & ~w2624;
assign w3259 = pi091 & ~pi115;
assign w3260 = pi092 & ~pi116;
assign w3261 = ~pi092 & pi116;
assign w3262 = pi094 & ~pi118;
assign w3263 = pi093 & ~pi117;
assign w3264 = ~w3262 & ~w3263;
assign w3265 = ~pi093 & pi117;
assign w3266 = ~w3261 & ~w3265;
assign w3267 = ~w3264 & w3266;
assign w3268 = ~w3259 & ~w3260;
assign w3269 = ~w3267 & w3268;
assign w3270 = ~pi091 & pi115;
assign w3271 = ~pi090 & pi114;
assign w3272 = ~w3270 & ~w3271;
assign w3273 = ~w3269 & w3272;
assign w3274 = pi090 & ~pi114;
assign w3275 = pi089 & ~pi113;
assign w3276 = ~w3274 & ~w3275;
assign w3277 = ~w3273 & w3276;
assign w3278 = ~pi089 & pi113;
assign w3279 = ~pi088 & pi112;
assign w3280 = ~w3278 & ~w3279;
assign w3281 = ~w3277 & w3280;
assign w3282 = pi088 & ~pi112;
assign w3283 = pi087 & ~pi111;
assign w3284 = ~w3282 & ~w3283;
assign w3285 = ~w3281 & w3284;
assign w3286 = ~pi087 & pi111;
assign w3287 = ~w3285 & ~w3286;
assign w3288 = ~w3258 & ~w3287;
assign w3289 = w2552 & w3288;
assign w3290 = w3257 & w3289;
assign w3291 = w2755 & w3290;
assign w3292 = w3054 & w3291;
assign w3293 = ~w2638 & w3292;
assign w3294 = ~w2637 & w3293;
assign w3295 = ~w342 & w2634;
assign w3296 = w3294 & ~w3295;
assign w3297 = pi007 & w3296;
assign w3298 = w1767 & ~w2570;
assign w3299 = w2534 & ~w2552;
assign w3300 = w2504 & ~w3299;
assign w3301 = w2582 & w3300;
assign w3302 = ~w3298 & w3301;
assign w3303 = ~w1230 & ~w2561;
assign w3304 = (w2387 & ~w2538) | (w2387 & w16232) | (~w2538 & w16232);
assign w3305 = ~w3303 & w3304;
assign w3306 = w3302 & w3305;
assign w3307 = pi005 & w3306;
assign w3308 = w1230 & ~w2538;
assign w3309 = w2582 & ~w3308;
assign w3310 = w1670 & w1728;
assign w3311 = (w3310 & ~w1423) | (w3310 & w16233) | (~w1423 & w16233);
assign w3312 = ~w467 & ~w2568;
assign w3313 = (w1199 & ~w2547) | (w1199 & w16234) | (~w2547 & w16234);
assign w3314 = w1106 & w1359;
assign w3315 = w1293 & w1418;
assign w3316 = w3314 & w3315;
assign w3317 = w1013 & ~w3313;
assign w3318 = w3316 & w3317;
assign w3319 = ~w3312 & w3318;
assign w3320 = w3311 & w3319;
assign w3321 = w1169 & ~w1755;
assign w3322 = ~w2561 & w3321;
assign w3323 = w3320 & w3322;
assign w3324 = w3309 & w3323;
assign w3325 = pi003 & w3324;
assign w3326 = ~w373 & ~w2552;
assign w3327 = w280 & w343;
assign w3328 = ~w3326 & w3327;
assign w3329 = (w3328 & w2561) | (w3328 & w16235) | (w2561 & w16235);
assign w3330 = w2634 & w3329;
assign w3331 = w404 & ~w1230;
assign w3332 = (w3331 & ~w1423) | (w3331 & w16236) | (~w1423 & w16236);
assign w3333 = (w404 & ~w2387) | (w404 & w16237) | (~w2387 & w16237);
assign w3334 = ~w3332 & ~w3333;
assign w3335 = w2582 & w3334;
assign w3336 = w917 & w3335;
assign w3337 = w3330 & w3336;
assign w3338 = pi001 & w3337;
assign w3339 = ~w2633 & ~w2636;
assign w3340 = ~w3325 & w3339;
assign w3341 = ~w3297 & ~w3307;
assign w3342 = ~w3338 & w3341;
assign w3343 = ~w2591 & w3340;
assign w3344 = w3342 & w3343;
assign w3345 = w2586 & ~w3306;
assign w3346 = (~w2582 & w2634) | (~w2582 & w17000) | (w2634 & w17000);
assign w3347 = w2587 & ~w3324;
assign w3348 = (~w3346 & w3324) | (~w3346 & w17001) | (w3324 & w17001);
assign w3349 = ~w3345 & w3348;
assign w3350 = w2634 & ~w3337;
assign w3351 = ~w3337 & w17002;
assign w3352 = w3349 & ~w3351;
assign w3353 = ~w2589 & w3352;
assign w3354 = pi006 & w3353;
assign w3355 = pi003 & w3321;
assign w3356 = w3312 & ~w3337;
assign w3357 = (~w1012 & ~w3294) | (~w1012 & w16238) | (~w3294 & w16238);
assign w3358 = ~w3356 & ~w3357;
assign w3359 = ~w3306 & w3308;
assign w3360 = w984 & ~w2631;
assign w3361 = (w3313 & ~w2585) | (w3313 & w17003) | (~w2585 & w17003);
assign w3362 = ~w3324 & ~w3346;
assign w3363 = w3310 & w3316;
assign w3364 = ~w3360 & w3363;
assign w3365 = ~w2561 & w3364;
assign w3366 = (w3365 & w3306) | (w3365 & w17004) | (w3306 & w17004);
assign w3367 = ~w3361 & w3362;
assign w3368 = w3366 & w3367;
assign w3369 = w3358 & w3368;
assign w3370 = w3355 & w3369;
assign w3371 = ~w2589 & w3299;
assign w3372 = (w2383 & ~w3294) | (w2383 & w16239) | (~w3294 & w16239);
assign w3373 = ~w3337 & w17005;
assign w3374 = ~w3371 & ~w3372;
assign w3375 = ~w3373 & w3374;
assign w3376 = ~w3306 & ~w3346;
assign w3377 = w3303 & ~w3324;
assign w3378 = (w1920 & ~w2538) | (w1920 & w16240) | (~w2538 & w16240);
assign w3379 = w2167 & w3378;
assign w3380 = ~w2354 & ~w2632;
assign w3381 = w2325 & w2504;
assign w3382 = ~w3380 & w3381;
assign w3383 = w3379 & w3382;
assign w3384 = ~w3377 & w3383;
assign w3385 = w3376 & w3384;
assign w3386 = w3384 & w16241;
assign w3387 = w3375 & w3386;
assign w3388 = pi005 & w3387;
assign w3389 = ~w3337 & w3295;
assign w3390 = (w3054 & ~w3294) | (w3054 & w16242) | (~w3294 & w16242);
assign w3391 = ~w2561 & ~w3324;
assign w3392 = ~w3324 & w2638;
assign w3393 = ~w2632 & w3258;
assign w3394 = w2637 & ~w3306;
assign w3395 = w2755 & ~w3393;
assign w3396 = w2589 & w3395;
assign w3397 = w3390 & w3396;
assign w3398 = ~w3392 & ~w3394;
assign w3399 = w3397 & w3398;
assign w3400 = w3257 & ~w3287;
assign w3401 = (w3400 & w3337) | (w3400 & w17533) | (w3337 & w17533);
assign w3402 = w3399 & w3401;
assign w3403 = pi007 & w3402;
assign w3404 = w2582 & ~w3337;
assign w3405 = ~w3337 & w17006;
assign w3406 = ~w3306 & ~w3334;
assign w3407 = ~w3324 & w16243;
assign w3408 = (w342 & ~w3293) | (w342 & w16244) | (~w3293 & w16244);
assign w3409 = w311 & ~w2632;
assign w3410 = w757 & w914;
assign w3411 = ~w2589 & w3326;
assign w3412 = w280 & w822;
assign w3413 = w3410 & w3412;
assign w3414 = ~w3409 & w3413;
assign w3415 = w2634 & w3414;
assign w3416 = ~w3408 & w3415;
assign w3417 = ~w3406 & w3416;
assign w3418 = ~w3407 & ~w3411;
assign w3419 = w3417 & w3418;
assign w3420 = w3405 & w3419;
assign w3421 = pi001 & w3420;
assign w3422 = pi104 & ~pi224;
assign w3423 = pi103 & ~pi223;
assign w3424 = ~pi104 & pi224;
assign w3425 = ~pi105 & pi225;
assign w3426 = pi106 & ~pi226;
assign w3427 = pi105 & ~pi225;
assign w3428 = pi107 & ~pi227;
assign w3429 = pi108 & ~pi228;
assign w3430 = pi109 & ~pi229;
assign w3431 = pi110 & ~pi230;
assign w3432 = ~w3430 & ~w3431;
assign w3433 = ~pi109 & pi229;
assign w3434 = ~pi108 & pi228;
assign w3435 = ~w3433 & ~w3434;
assign w3436 = ~w3432 & w3435;
assign w3437 = ~w3428 & ~w3429;
assign w3438 = ~pi106 & pi226;
assign w3439 = ~pi107 & pi227;
assign w3440 = ~w3438 & ~w3439;
assign w3441 = (w3440 & w3436) | (w3440 & w17534) | (w3436 & w17534);
assign w3442 = ~w3426 & ~w3427;
assign w3443 = ~w3441 & w3442;
assign w3444 = ~w3424 & ~w3425;
assign w3445 = ~w3443 & w3444;
assign w3446 = ~w3422 & ~w3423;
assign w3447 = ~w3445 & w3446;
assign w3448 = ~pi103 & pi223;
assign w3449 = ~w3447 & ~w3448;
assign w3450 = pi104 & ~pi216;
assign w3451 = pi103 & ~pi215;
assign w3452 = ~pi104 & pi216;
assign w3453 = ~pi105 & pi217;
assign w3454 = pi106 & ~pi218;
assign w3455 = pi105 & ~pi217;
assign w3456 = pi107 & ~pi219;
assign w3457 = pi108 & ~pi220;
assign w3458 = pi109 & ~pi221;
assign w3459 = pi110 & ~pi222;
assign w3460 = ~w3458 & ~w3459;
assign w3461 = ~pi109 & pi221;
assign w3462 = ~pi108 & pi220;
assign w3463 = ~w3461 & ~w3462;
assign w3464 = ~w3460 & w3463;
assign w3465 = ~w3456 & ~w3457;
assign w3466 = ~pi106 & pi218;
assign w3467 = ~pi107 & pi219;
assign w3468 = ~w3466 & ~w3467;
assign w3469 = (w3468 & w3464) | (w3468 & w17535) | (w3464 & w17535);
assign w3470 = ~w3454 & ~w3455;
assign w3471 = ~w3469 & w3470;
assign w3472 = ~w3452 & ~w3453;
assign w3473 = ~w3471 & w3472;
assign w3474 = ~w3450 & ~w3451;
assign w3475 = ~w3473 & w3474;
assign w3476 = ~pi103 & pi215;
assign w3477 = ~w3475 & ~w3476;
assign w3478 = ~w3449 & ~w3477;
assign w3479 = pi104 & ~pi200;
assign w3480 = pi103 & ~pi199;
assign w3481 = ~pi104 & pi200;
assign w3482 = ~pi105 & pi201;
assign w3483 = pi105 & ~pi201;
assign w3484 = pi106 & ~pi202;
assign w3485 = ~pi106 & pi202;
assign w3486 = ~pi107 & pi203;
assign w3487 = pi108 & ~pi204;
assign w3488 = pi107 & ~pi203;
assign w3489 = pi109 & ~pi205;
assign w3490 = pi110 & ~pi206;
assign w3491 = ~w3489 & ~w3490;
assign w3492 = ~pi109 & pi205;
assign w3493 = ~pi108 & pi204;
assign w3494 = ~w3492 & ~w3493;
assign w3495 = ~w3491 & w3494;
assign w3496 = ~w3487 & ~w3488;
assign w3497 = ~w3485 & ~w3486;
assign w3498 = (w3497 & w3495) | (w3497 & w17536) | (w3495 & w17536);
assign w3499 = ~w3483 & ~w3484;
assign w3500 = ~w3498 & w3499;
assign w3501 = ~w3481 & ~w3482;
assign w3502 = ~w3500 & w3501;
assign w3503 = ~w3479 & ~w3480;
assign w3504 = ~w3502 & w3503;
assign w3505 = ~pi103 & pi199;
assign w3506 = ~w3504 & ~w3505;
assign w3507 = pi104 & ~pi208;
assign w3508 = pi103 & ~pi207;
assign w3509 = ~pi104 & pi208;
assign w3510 = ~pi105 & pi209;
assign w3511 = pi106 & ~pi210;
assign w3512 = pi105 & ~pi209;
assign w3513 = pi107 & ~pi211;
assign w3514 = pi108 & ~pi212;
assign w3515 = pi109 & ~pi213;
assign w3516 = pi110 & ~pi214;
assign w3517 = ~w3515 & ~w3516;
assign w3518 = ~pi109 & pi213;
assign w3519 = ~pi108 & pi212;
assign w3520 = ~w3518 & ~w3519;
assign w3521 = ~w3517 & w3520;
assign w3522 = ~w3513 & ~w3514;
assign w3523 = ~pi106 & pi210;
assign w3524 = ~pi107 & pi211;
assign w3525 = ~w3523 & ~w3524;
assign w3526 = (w3525 & w3521) | (w3525 & w17537) | (w3521 & w17537);
assign w3527 = ~w3511 & ~w3512;
assign w3528 = ~w3526 & w3527;
assign w3529 = ~w3509 & ~w3510;
assign w3530 = ~w3528 & w3529;
assign w3531 = ~w3507 & ~w3508;
assign w3532 = ~w3530 & w3531;
assign w3533 = ~pi103 & pi207;
assign w3534 = ~w3532 & ~w3533;
assign w3535 = ~w3506 & ~w3534;
assign w3536 = w3478 & w3535;
assign w3537 = pi103 & ~pi191;
assign w3538 = ~pi103 & pi191;
assign w3539 = pi104 & ~pi192;
assign w3540 = ~pi104 & pi192;
assign w3541 = ~pi105 & pi193;
assign w3542 = pi105 & ~pi193;
assign w3543 = pi106 & ~pi194;
assign w3544 = pi107 & ~pi195;
assign w3545 = pi108 & ~pi196;
assign w3546 = ~pi108 & pi196;
assign w3547 = pi109 & ~pi197;
assign w3548 = pi110 & ~pi198;
assign w3549 = ~w3547 & ~w3548;
assign w3550 = ~pi109 & pi197;
assign w3551 = ~w3546 & ~w3550;
assign w3552 = ~w3549 & w3551;
assign w3553 = ~w3544 & ~w3545;
assign w3554 = ~w3552 & w3553;
assign w3555 = ~pi106 & pi194;
assign w3556 = ~pi107 & pi195;
assign w3557 = ~w3555 & ~w3556;
assign w3558 = ~w3554 & w3557;
assign w3559 = ~w3542 & ~w3543;
assign w3560 = ~w3558 & w3559;
assign w3561 = ~w3540 & ~w3541;
assign w3562 = ~w3560 & w3561;
assign w3563 = ~w3539 & ~w3562;
assign w3564 = ~w3538 & ~w3563;
assign w3565 = ~w3537 & ~w3564;
assign w3566 = w3536 & w3565;
assign w3567 = ~pi103 & pi167;
assign w3568 = pi103 & ~pi167;
assign w3569 = pi104 & ~pi168;
assign w3570 = pi105 & ~pi169;
assign w3571 = pi106 & ~pi170;
assign w3572 = ~pi106 & pi170;
assign w3573 = ~pi107 & pi171;
assign w3574 = pi107 & ~pi171;
assign w3575 = pi108 & ~pi172;
assign w3576 = ~pi109 & pi173;
assign w3577 = pi109 & ~pi173;
assign w3578 = pi110 & ~pi174;
assign w3579 = ~w3577 & ~w3578;
assign w3580 = ~pi108 & pi172;
assign w3581 = ~w3576 & ~w3580;
assign w3582 = ~w3579 & w3581;
assign w3583 = ~w3574 & ~w3575;
assign w3584 = ~w3582 & w3583;
assign w3585 = ~w3572 & ~w3573;
assign w3586 = ~w3584 & w3585;
assign w3587 = ~w3570 & ~w3571;
assign w3588 = ~w3586 & w3587;
assign w3589 = ~pi104 & pi168;
assign w3590 = ~pi105 & pi169;
assign w3591 = ~w3589 & ~w3590;
assign w3592 = ~w3588 & w3591;
assign w3593 = ~w3568 & ~w3569;
assign w3594 = ~w3592 & w3593;
assign w3595 = ~w3567 & ~w3594;
assign w3596 = ~pi103 & pi175;
assign w3597 = ~pi104 & pi176;
assign w3598 = ~pi105 & pi177;
assign w3599 = pi106 & ~pi178;
assign w3600 = pi105 & ~pi177;
assign w3601 = ~pi106 & pi178;
assign w3602 = ~pi107 & pi179;
assign w3603 = pi109 & ~pi181;
assign w3604 = ~pi109 & pi181;
assign w3605 = pi110 & ~pi182;
assign w3606 = ~w3604 & w3605;
assign w3607 = (~pi180 & w3606) | (~pi180 & w17538) | (w3606 & w17538);
assign w3608 = pi107 & ~pi179;
assign w3609 = ~w3606 & w17539;
assign w3610 = pi108 & ~w3609;
assign w3611 = ~w3607 & ~w3608;
assign w3612 = ~w3610 & w3611;
assign w3613 = ~w3601 & ~w3602;
assign w3614 = ~w3612 & w3613;
assign w3615 = ~w3599 & ~w3600;
assign w3616 = ~w3614 & w3615;
assign w3617 = ~w3597 & ~w3598;
assign w3618 = ~w3616 & w3617;
assign w3619 = pi103 & ~pi175;
assign w3620 = pi104 & ~pi176;
assign w3621 = ~w3619 & ~w3620;
assign w3622 = ~w3618 & w3621;
assign w3623 = ~w3596 & ~w3622;
assign w3624 = ~w3595 & ~w3623;
assign w3625 = w3566 & w3624;
assign w3626 = ~pi103 & pi151;
assign w3627 = ~pi104 & pi152;
assign w3628 = ~pi105 & pi153;
assign w3629 = pi105 & ~pi153;
assign w3630 = pi106 & ~pi154;
assign w3631 = ~pi107 & pi155;
assign w3632 = ~pi106 & pi154;
assign w3633 = pi109 & ~pi157;
assign w3634 = ~pi109 & pi157;
assign w3635 = pi110 & ~pi158;
assign w3636 = ~w3634 & w3635;
assign w3637 = ~w3633 & ~w3636;
assign w3638 = ~pi156 & ~w3637;
assign w3639 = pi107 & ~pi155;
assign w3640 = pi156 & w3637;
assign w3641 = pi108 & ~w3640;
assign w3642 = ~w3638 & ~w3639;
assign w3643 = ~w3641 & w3642;
assign w3644 = ~w3631 & ~w3632;
assign w3645 = ~w3643 & w3644;
assign w3646 = ~w3629 & ~w3630;
assign w3647 = ~w3645 & w3646;
assign w3648 = ~w3627 & ~w3628;
assign w3649 = ~w3647 & w3648;
assign w3650 = pi103 & ~pi151;
assign w3651 = pi104 & ~pi152;
assign w3652 = ~w3650 & ~w3651;
assign w3653 = ~w3649 & w3652;
assign w3654 = ~w3626 & ~w3653;
assign w3655 = ~pi103 & pi159;
assign w3656 = ~pi104 & pi160;
assign w3657 = ~pi105 & pi161;
assign w3658 = pi105 & ~pi161;
assign w3659 = pi106 & ~pi162;
assign w3660 = ~pi106 & pi162;
assign w3661 = ~pi107 & pi163;
assign w3662 = pi109 & ~pi165;
assign w3663 = ~pi109 & pi165;
assign w3664 = pi110 & ~pi166;
assign w3665 = ~w3663 & w3664;
assign w3666 = ~w3662 & ~w3665;
assign w3667 = ~pi164 & ~w3666;
assign w3668 = pi107 & ~pi163;
assign w3669 = pi164 & w3666;
assign w3670 = pi108 & ~w3669;
assign w3671 = ~w3667 & ~w3668;
assign w3672 = ~w3670 & w3671;
assign w3673 = ~w3660 & ~w3661;
assign w3674 = ~w3672 & w3673;
assign w3675 = ~w3658 & ~w3659;
assign w3676 = ~w3674 & w3675;
assign w3677 = ~w3656 & ~w3657;
assign w3678 = ~w3676 & w3677;
assign w3679 = pi103 & ~pi159;
assign w3680 = pi104 & ~pi160;
assign w3681 = ~w3679 & ~w3680;
assign w3682 = ~w3678 & w3681;
assign w3683 = ~w3655 & ~w3682;
assign w3684 = ~w3654 & ~w3683;
assign w3685 = w3625 & w3684;
assign w3686 = ~pi103 & pi135;
assign w3687 = pi103 & ~pi135;
assign w3688 = pi104 & ~pi136;
assign w3689 = ~pi104 & pi136;
assign w3690 = ~pi105 & pi137;
assign w3691 = pi105 & ~pi137;
assign w3692 = pi106 & ~pi138;
assign w3693 = pi107 & ~pi139;
assign w3694 = pi108 & ~pi140;
assign w3695 = ~pi109 & pi141;
assign w3696 = pi109 & ~pi141;
assign w3697 = pi110 & ~pi142;
assign w3698 = ~w3696 & ~w3697;
assign w3699 = ~pi108 & pi140;
assign w3700 = ~w3695 & ~w3699;
assign w3701 = ~w3698 & w3700;
assign w3702 = ~w3693 & ~w3694;
assign w3703 = ~w3701 & w3702;
assign w3704 = ~pi106 & pi138;
assign w3705 = ~pi107 & pi139;
assign w3706 = ~w3704 & ~w3705;
assign w3707 = ~w3703 & w3706;
assign w3708 = ~w3691 & ~w3692;
assign w3709 = ~w3707 & w3708;
assign w3710 = ~w3689 & ~w3690;
assign w3711 = ~w3709 & w3710;
assign w3712 = ~w3687 & ~w3688;
assign w3713 = ~w3711 & w3712;
assign w3714 = ~w3686 & ~w3713;
assign w3715 = ~pi103 & pi143;
assign w3716 = pi104 & ~pi144;
assign w3717 = pi103 & ~pi143;
assign w3718 = ~pi105 & pi145;
assign w3719 = ~pi104 & pi144;
assign w3720 = pi105 & ~pi145;
assign w3721 = pi106 & ~pi146;
assign w3722 = ~pi107 & pi147;
assign w3723 = ~pi106 & pi146;
assign w3724 = pi109 & ~pi149;
assign w3725 = ~pi109 & pi149;
assign w3726 = pi110 & ~pi150;
assign w3727 = ~w3725 & w3726;
assign w3728 = ~w3724 & ~w3727;
assign w3729 = ~pi148 & ~w3728;
assign w3730 = pi107 & ~pi147;
assign w3731 = pi148 & w3728;
assign w3732 = pi108 & ~w3731;
assign w3733 = ~w3729 & ~w3730;
assign w3734 = ~w3732 & w3733;
assign w3735 = ~w3722 & ~w3723;
assign w3736 = ~w3734 & w3735;
assign w3737 = ~w3720 & ~w3721;
assign w3738 = ~w3736 & w3737;
assign w3739 = ~w3718 & ~w3719;
assign w3740 = ~w3738 & w3739;
assign w3741 = ~w3716 & ~w3717;
assign w3742 = ~w3740 & w3741;
assign w3743 = ~w3715 & ~w3742;
assign w3744 = ~w3714 & ~w3743;
assign w3745 = w3685 & w3744;
assign w3746 = ~pi104 & pi256;
assign w3747 = ~pi105 & pi257;
assign w3748 = pi105 & ~pi257;
assign w3749 = pi106 & ~pi258;
assign w3750 = ~pi106 & pi258;
assign w3751 = ~pi107 & pi259;
assign w3752 = pi109 & ~pi261;
assign w3753 = ~pi109 & pi261;
assign w3754 = pi110 & ~pi262;
assign w3755 = ~w3753 & w3754;
assign w3756 = (~pi260 & w3755) | (~pi260 & w17540) | (w3755 & w17540);
assign w3757 = pi107 & ~pi259;
assign w3758 = ~w3755 & w17541;
assign w3759 = pi108 & ~w3758;
assign w3760 = ~w3756 & ~w3757;
assign w3761 = ~w3759 & w3760;
assign w3762 = ~w3750 & ~w3751;
assign w3763 = ~w3761 & w3762;
assign w3764 = ~w3748 & ~w3749;
assign w3765 = ~w3763 & w3764;
assign w3766 = ~w3746 & ~w3747;
assign w3767 = ~w3765 & w3766;
assign w3768 = pi103 & ~pi255;
assign w3769 = pi104 & ~pi256;
assign w3770 = ~w3768 & ~w3769;
assign w3771 = ~w3767 & w3770;
assign w3772 = ~pi103 & pi255;
assign w3773 = ~w3771 & ~w3772;
assign w3774 = ~pi105 & pi241;
assign w3775 = ~pi104 & pi240;
assign w3776 = pi106 & ~pi242;
assign w3777 = pi105 & ~pi241;
assign w3778 = ~pi106 & pi242;
assign w3779 = ~pi107 & pi243;
assign w3780 = pi108 & ~pi244;
assign w3781 = pi107 & ~pi243;
assign w3782 = ~pi108 & pi244;
assign w3783 = pi109 & ~pi245;
assign w3784 = ~pi109 & pi245;
assign w3785 = pi110 & ~pi246;
assign w3786 = ~w3784 & w3785;
assign w3787 = (~w3782 & w3786) | (~w3782 & w17542) | (w3786 & w17542);
assign w3788 = ~w3780 & ~w3781;
assign w3789 = ~w3787 & w3788;
assign w3790 = ~w3778 & ~w3779;
assign w3791 = ~w3789 & w3790;
assign w3792 = ~w3776 & ~w3777;
assign w3793 = ~w3791 & w3792;
assign w3794 = ~w3774 & ~w3775;
assign w3795 = ~w3793 & w3794;
assign w3796 = pi104 & ~pi240;
assign w3797 = pi103 & ~pi239;
assign w3798 = ~w3796 & ~w3797;
assign w3799 = ~w3795 & w3798;
assign w3800 = ~pi103 & pi239;
assign w3801 = ~w3799 & ~w3800;
assign w3802 = ~pi103 & pi231;
assign w3803 = pi103 & ~pi231;
assign w3804 = pi104 & ~pi232;
assign w3805 = pi105 & ~pi233;
assign w3806 = pi106 & ~pi234;
assign w3807 = ~pi106 & pi234;
assign w3808 = ~pi107 & pi235;
assign w3809 = ~pi108 & pi236;
assign w3810 = pi109 & ~pi237;
assign w3811 = pi110 & ~pi238;
assign w3812 = ~w3810 & ~w3811;
assign w3813 = ~pi109 & pi237;
assign w3814 = ~w3809 & ~w3813;
assign w3815 = ~w3812 & w3814;
assign w3816 = pi107 & ~pi235;
assign w3817 = pi108 & ~pi236;
assign w3818 = ~w3816 & ~w3817;
assign w3819 = ~w3815 & w3818;
assign w3820 = ~w3807 & ~w3808;
assign w3821 = ~w3819 & w3820;
assign w3822 = ~w3805 & ~w3806;
assign w3823 = ~w3821 & w3822;
assign w3824 = ~pi104 & pi232;
assign w3825 = ~pi105 & pi233;
assign w3826 = ~w3824 & ~w3825;
assign w3827 = ~w3823 & w3826;
assign w3828 = ~w3803 & ~w3804;
assign w3829 = ~w3827 & w3828;
assign w3830 = ~w3802 & ~w3829;
assign w3831 = ~w3801 & ~w3830;
assign w3832 = ~w3773 & w3831;
assign w3833 = ~pi104 & pi248;
assign w3834 = ~pi105 & pi249;
assign w3835 = pi106 & ~pi250;
assign w3836 = pi105 & ~pi249;
assign w3837 = ~pi106 & pi250;
assign w3838 = ~pi107 & pi251;
assign w3839 = pi109 & ~pi253;
assign w3840 = ~pi109 & pi253;
assign w3841 = pi110 & ~pi254;
assign w3842 = ~w3840 & w3841;
assign w3843 = (~pi252 & w3842) | (~pi252 & w17543) | (w3842 & w17543);
assign w3844 = pi107 & ~pi251;
assign w3845 = ~w3842 & w17544;
assign w3846 = pi108 & ~w3845;
assign w3847 = ~w3843 & ~w3844;
assign w3848 = ~w3846 & w3847;
assign w3849 = ~w3837 & ~w3838;
assign w3850 = ~w3848 & w3849;
assign w3851 = ~w3835 & ~w3836;
assign w3852 = ~w3850 & w3851;
assign w3853 = ~w3833 & ~w3834;
assign w3854 = ~w3852 & w3853;
assign w3855 = pi103 & ~pi247;
assign w3856 = pi104 & ~pi248;
assign w3857 = ~w3855 & ~w3856;
assign w3858 = ~w3854 & w3857;
assign w3859 = ~pi103 & pi247;
assign w3860 = ~w3858 & ~w3859;
assign w3861 = ~pi104 & pi272;
assign w3862 = ~pi105 & pi273;
assign w3863 = pi106 & ~pi274;
assign w3864 = pi105 & ~pi273;
assign w3865 = ~pi106 & pi274;
assign w3866 = ~pi107 & pi275;
assign w3867 = pi108 & ~pi276;
assign w3868 = pi107 & ~pi275;
assign w3869 = ~pi108 & pi276;
assign w3870 = pi109 & ~pi277;
assign w3871 = ~pi109 & pi277;
assign w3872 = pi110 & ~pi278;
assign w3873 = ~w3871 & w3872;
assign w3874 = (~w3869 & w3873) | (~w3869 & w17545) | (w3873 & w17545);
assign w3875 = ~w3867 & ~w3868;
assign w3876 = ~w3874 & w3875;
assign w3877 = ~w3865 & ~w3866;
assign w3878 = ~w3876 & w3877;
assign w3879 = ~w3863 & ~w3864;
assign w3880 = ~w3878 & w3879;
assign w3881 = ~w3861 & ~w3862;
assign w3882 = ~w3880 & w3881;
assign w3883 = pi104 & ~pi272;
assign w3884 = pi103 & ~pi271;
assign w3885 = ~w3883 & ~w3884;
assign w3886 = ~w3882 & w3885;
assign w3887 = ~pi103 & pi271;
assign w3888 = ~w3886 & ~w3887;
assign w3889 = ~pi103 & pi263;
assign w3890 = pi103 & ~pi263;
assign w3891 = pi104 & ~pi264;
assign w3892 = pi105 & ~pi265;
assign w3893 = pi106 & ~pi266;
assign w3894 = ~pi106 & pi266;
assign w3895 = ~pi107 & pi267;
assign w3896 = ~pi108 & pi268;
assign w3897 = pi109 & ~pi269;
assign w3898 = pi110 & ~pi270;
assign w3899 = ~w3897 & ~w3898;
assign w3900 = ~pi109 & pi269;
assign w3901 = ~w3896 & ~w3900;
assign w3902 = ~w3899 & w3901;
assign w3903 = pi107 & ~pi267;
assign w3904 = pi108 & ~pi268;
assign w3905 = ~w3903 & ~w3904;
assign w3906 = ~w3902 & w3905;
assign w3907 = ~w3894 & ~w3895;
assign w3908 = ~w3906 & w3907;
assign w3909 = ~w3892 & ~w3893;
assign w3910 = ~w3908 & w3909;
assign w3911 = ~pi104 & pi264;
assign w3912 = ~pi105 & pi265;
assign w3913 = ~w3911 & ~w3912;
assign w3914 = ~w3910 & w3913;
assign w3915 = ~w3890 & ~w3891;
assign w3916 = ~w3914 & w3915;
assign w3917 = ~w3889 & ~w3916;
assign w3918 = ~w3888 & ~w3917;
assign w3919 = ~w3860 & w3918;
assign w3920 = w3832 & w3919;
assign w3921 = ~pi103 & pi183;
assign w3922 = pi104 & ~pi184;
assign w3923 = pi103 & ~pi183;
assign w3924 = pi105 & ~pi185;
assign w3925 = pi106 & ~pi186;
assign w3926 = ~pi106 & pi186;
assign w3927 = ~pi107 & pi187;
assign w3928 = pi107 & ~pi187;
assign w3929 = pi108 & ~pi188;
assign w3930 = ~pi109 & pi189;
assign w3931 = pi109 & ~pi189;
assign w3932 = pi110 & ~pi190;
assign w3933 = ~w3931 & ~w3932;
assign w3934 = ~pi108 & pi188;
assign w3935 = ~w3930 & ~w3934;
assign w3936 = ~w3933 & w3935;
assign w3937 = ~w3928 & ~w3929;
assign w3938 = ~w3936 & w3937;
assign w3939 = ~w3926 & ~w3927;
assign w3940 = ~w3938 & w3939;
assign w3941 = ~w3924 & ~w3925;
assign w3942 = ~w3940 & w3941;
assign w3943 = ~pi104 & pi184;
assign w3944 = ~pi105 & pi185;
assign w3945 = ~w3943 & ~w3944;
assign w3946 = ~w3942 & w3945;
assign w3947 = ~w3922 & ~w3923;
assign w3948 = ~w3946 & w3947;
assign w3949 = ~w3921 & ~w3948;
assign w3950 = ~pi103 & pi127;
assign w3951 = pi104 & ~pi128;
assign w3952 = pi103 & ~pi127;
assign w3953 = ~pi104 & pi128;
assign w3954 = ~pi105 & pi129;
assign w3955 = pi106 & ~pi130;
assign w3956 = pi105 & ~pi129;
assign w3957 = pi107 & ~pi131;
assign w3958 = pi108 & ~pi132;
assign w3959 = ~pi109 & pi133;
assign w3960 = pi109 & ~pi133;
assign w3961 = pi110 & ~pi134;
assign w3962 = ~w3960 & ~w3961;
assign w3963 = ~pi108 & pi132;
assign w3964 = ~w3959 & ~w3963;
assign w3965 = ~w3962 & w3964;
assign w3966 = ~w3957 & ~w3958;
assign w3967 = ~w3965 & w3966;
assign w3968 = ~pi106 & pi130;
assign w3969 = ~pi107 & pi131;
assign w3970 = ~w3968 & ~w3969;
assign w3971 = ~w3967 & w3970;
assign w3972 = ~w3955 & ~w3956;
assign w3973 = ~w3971 & w3972;
assign w3974 = ~w3953 & ~w3954;
assign w3975 = ~w3973 & w3974;
assign w3976 = ~w3951 & ~w3952;
assign w3977 = ~w3975 & w3976;
assign w3978 = ~w3950 & ~w3977;
assign w3979 = ~w3949 & ~w3978;
assign w3980 = w3920 & w3979;
assign w3981 = ~pi103 & pi119;
assign w3982 = pi103 & ~pi119;
assign w3983 = pi104 & ~pi120;
assign w3984 = ~pi104 & pi120;
assign w3985 = ~pi105 & pi121;
assign w3986 = pi105 & ~pi121;
assign w3987 = pi106 & ~pi122;
assign w3988 = ~pi107 & pi123;
assign w3989 = ~pi106 & pi122;
assign w3990 = pi107 & ~pi123;
assign w3991 = pi108 & ~pi124;
assign w3992 = ~pi108 & pi124;
assign w3993 = pi109 & ~pi125;
assign w3994 = ~pi109 & pi125;
assign w3995 = pi110 & ~pi126;
assign w3996 = ~w3994 & w3995;
assign w3997 = ~w3993 & ~w3996;
assign w3998 = ~w3992 & ~w3997;
assign w3999 = ~w3990 & ~w3991;
assign w4000 = ~w3998 & w3999;
assign w4001 = ~w3988 & ~w3989;
assign w4002 = ~w4000 & w4001;
assign w4003 = ~w3986 & ~w3987;
assign w4004 = ~w4002 & w4003;
assign w4005 = ~w3984 & ~w3985;
assign w4006 = ~w4004 & w4005;
assign w4007 = ~w3982 & ~w3983;
assign w4008 = ~w4006 & w4007;
assign w4009 = ~w3981 & ~w4008;
assign w4010 = ~pi104 & pi112;
assign w4011 = ~pi105 & pi113;
assign w4012 = pi105 & ~pi113;
assign w4013 = pi106 & ~pi114;
assign w4014 = ~pi106 & pi114;
assign w4015 = ~pi107 & pi115;
assign w4016 = pi109 & ~pi117;
assign w4017 = ~pi109 & pi117;
assign w4018 = pi110 & ~pi118;
assign w4019 = ~w4017 & w4018;
assign w4020 = ~w4016 & ~w4019;
assign w4021 = ~pi116 & ~w4020;
assign w4022 = pi107 & ~pi115;
assign w4023 = pi116 & w4020;
assign w4024 = pi108 & ~w4023;
assign w4025 = ~w4021 & ~w4022;
assign w4026 = ~w4024 & w4025;
assign w4027 = ~w4014 & ~w4015;
assign w4028 = ~w4026 & w4027;
assign w4029 = ~w4012 & ~w4013;
assign w4030 = ~w4028 & w4029;
assign w4031 = ~w4010 & ~w4011;
assign w4032 = ~w4030 & w4031;
assign w4033 = pi104 & ~pi112;
assign w4034 = pi103 & ~pi111;
assign w4035 = ~w4033 & ~w4034;
assign w4036 = ~w4032 & w4035;
assign w4037 = ~pi103 & pi111;
assign w4038 = ~w4036 & ~w4037;
assign w4039 = (~w2502 & ~w2538) | (~w2502 & w17546) | (~w2538 & w17546);
assign w4040 = ~w3306 & w4039;
assign w4041 = ~w3324 & w16245;
assign w4042 = ~w278 & w2634;
assign w4043 = ~w3337 & w4042;
assign w4044 = ~w2667 & ~w4009;
assign w4045 = ~w4038 & w4044;
assign w4046 = w2632 & w4045;
assign w4047 = w3980 & w4046;
assign w4048 = w3745 & w4047;
assign w4049 = (w4048 & w3306) | (w4048 & w17007) | (w3306 & w17007);
assign w4050 = ~w4041 & ~w4043;
assign w4051 = w4049 & w4050;
assign w4052 = pi009 & w4051;
assign w4053 = w717 & w720;
assign w4054 = w696 & ~w4053;
assign w4055 = ~w3286 & ~w4037;
assign w4056 = ~w2231 & w4055;
assign w4057 = w2596 & w4056;
assign w4058 = ~w1382 & w1385;
assign w4059 = w1363 & ~w4058;
assign w4060 = ~w983 & ~w4059;
assign w4061 = w2628 & w4060;
assign w4062 = ~w2259 & ~w3285;
assign w4063 = w2629 & w4062;
assign w4064 = ~w1360 & w2549;
assign w4065 = w4057 & w4064;
assign w4066 = ~w4054 & w4065;
assign w4067 = ~w4036 & w4066;
assign w4068 = w4063 & w4067;
assign w4069 = w4061 & w4068;
assign w4070 = w2548 & w4069;
assign w4071 = ~w693 & w4070;
assign w4072 = pi010 & w4071;
assign w4073 = ~w984 & w3391;
assign w4074 = ~w311 & w2634;
assign w4075 = ~w3337 & w4074;
assign w4076 = (~w3258 & ~w3294) | (~w3258 & w16246) | (~w3294 & w16246);
assign w4077 = w2354 & ~w2540;
assign w4078 = ~w3306 & w4077;
assign w4079 = w2589 & ~w2632;
assign w4080 = ~w4075 & w4079;
assign w4081 = ~w4076 & ~w4078;
assign w4082 = w4080 & w4081;
assign w4083 = ~w4073 & w4082;
assign w4084 = pi008 & w4083;
assign w4085 = ~w4052 & ~w4072;
assign w4086 = ~w3354 & w4085;
assign w4087 = ~w3370 & ~w3388;
assign w4088 = ~w3403 & ~w3421;
assign w4089 = ~w4084 & w4088;
assign w4090 = w4086 & w4087;
assign w4091 = w4089 & w4090;
assign w4092 = w3345 & ~w3387;
assign w4093 = w3321 & w3358;
assign w4094 = w3368 & w4093;
assign w4095 = w3347 & ~w4094;
assign w4096 = ~w4092 & ~w4095;
assign w4097 = ~w3346 & ~w3352;
assign w4098 = (w3351 & ~w3419) | (w3351 & w17547) | (~w3419 & w17547);
assign w4099 = w4097 & ~w4098;
assign w4100 = w4096 & w4099;
assign w4101 = pi006 & w4100;
assign w4102 = ~w2561 & ~w4094;
assign w4103 = ~w4094 & w3391;
assign w4104 = ~w4094 & w17548;
assign w4105 = (~w4009 & ~w4050) | (~w4009 & w17008) | (~w4050 & w17008);
assign w4106 = ~pi119 & pi135;
assign w4107 = pi119 & ~pi135;
assign w4108 = pi120 & ~pi136;
assign w4109 = ~pi121 & pi137;
assign w4110 = ~pi120 & pi136;
assign w4111 = pi121 & ~pi137;
assign w4112 = pi122 & ~pi138;
assign w4113 = ~pi122 & pi138;
assign w4114 = ~pi123 & pi139;
assign w4115 = pi125 & ~pi141;
assign w4116 = ~pi125 & pi141;
assign w4117 = pi126 & ~pi142;
assign w4118 = ~w4116 & w4117;
assign w4119 = ~w4115 & ~w4118;
assign w4120 = ~pi140 & ~w4119;
assign w4121 = pi123 & ~pi139;
assign w4122 = pi140 & w4119;
assign w4123 = pi124 & ~w4122;
assign w4124 = ~w4120 & ~w4121;
assign w4125 = ~w4123 & w4124;
assign w4126 = ~w4113 & ~w4114;
assign w4127 = ~w4125 & w4126;
assign w4128 = ~w4111 & ~w4112;
assign w4129 = ~w4127 & w4128;
assign w4130 = ~w4109 & ~w4110;
assign w4131 = ~w4129 & w4130;
assign w4132 = ~w4107 & ~w4108;
assign w4133 = ~w4131 & w4132;
assign w4134 = ~w4106 & ~w4133;
assign w4135 = ~pi119 & pi143;
assign w4136 = pi119 & ~pi143;
assign w4137 = ~pi120 & pi144;
assign w4138 = pi120 & ~pi144;
assign w4139 = ~pi121 & pi145;
assign w4140 = pi121 & ~pi145;
assign w4141 = pi122 & ~pi146;
assign w4142 = ~pi122 & pi146;
assign w4143 = ~pi123 & pi147;
assign w4144 = pi125 & ~pi149;
assign w4145 = ~pi125 & pi149;
assign w4146 = pi126 & ~pi150;
assign w4147 = ~w4145 & w4146;
assign w4148 = ~w4144 & ~w4147;
assign w4149 = ~pi148 & ~w4148;
assign w4150 = pi123 & ~pi147;
assign w4151 = pi148 & w4148;
assign w4152 = pi124 & ~w4151;
assign w4153 = ~w4149 & ~w4150;
assign w4154 = ~w4152 & w4153;
assign w4155 = ~w4142 & ~w4143;
assign w4156 = ~w4154 & w4155;
assign w4157 = ~w4140 & ~w4141;
assign w4158 = ~w4156 & w4157;
assign w4159 = ~w4139 & ~w4158;
assign w4160 = ~w4138 & ~w4159;
assign w4161 = ~w4137 & ~w4160;
assign w4162 = ~w4136 & ~w4161;
assign w4163 = ~w4135 & ~w4162;
assign w4164 = ~pi119 & pi255;
assign w4165 = pi120 & ~pi256;
assign w4166 = pi119 & ~pi255;
assign w4167 = ~pi120 & pi256;
assign w4168 = ~pi121 & pi257;
assign w4169 = pi121 & ~pi257;
assign w4170 = pi122 & ~pi258;
assign w4171 = ~pi122 & pi258;
assign w4172 = ~pi123 & pi259;
assign w4173 = pi123 & ~pi259;
assign w4174 = pi124 & ~pi260;
assign w4175 = ~pi125 & pi261;
assign w4176 = pi125 & ~pi261;
assign w4177 = pi126 & ~pi262;
assign w4178 = ~w4176 & ~w4177;
assign w4179 = ~pi124 & pi260;
assign w4180 = ~w4175 & ~w4179;
assign w4181 = ~w4178 & w4180;
assign w4182 = ~w4173 & ~w4174;
assign w4183 = ~w4181 & w4182;
assign w4184 = ~w4171 & ~w4172;
assign w4185 = ~w4183 & w4184;
assign w4186 = ~w4169 & ~w4170;
assign w4187 = ~w4185 & w4186;
assign w4188 = ~w4167 & ~w4168;
assign w4189 = ~w4187 & w4188;
assign w4190 = ~w4165 & ~w4166;
assign w4191 = ~w4189 & w4190;
assign w4192 = ~w4164 & ~w4191;
assign w4193 = ~pi119 & pi263;
assign w4194 = pi119 & ~pi263;
assign w4195 = pi120 & ~pi264;
assign w4196 = ~pi120 & pi264;
assign w4197 = ~pi121 & pi265;
assign w4198 = pi121 & ~pi265;
assign w4199 = pi122 & ~pi266;
assign w4200 = ~pi122 & pi266;
assign w4201 = ~pi123 & pi267;
assign w4202 = pi125 & ~pi269;
assign w4203 = ~pi125 & pi269;
assign w4204 = pi126 & ~pi270;
assign w4205 = ~w4203 & w4204;
assign w4206 = ~w4202 & ~w4205;
assign w4207 = ~pi268 & ~w4206;
assign w4208 = pi123 & ~pi267;
assign w4209 = pi268 & w4206;
assign w4210 = pi124 & ~w4209;
assign w4211 = ~w4207 & ~w4208;
assign w4212 = ~w4210 & w4211;
assign w4213 = ~w4200 & ~w4201;
assign w4214 = ~w4212 & w4213;
assign w4215 = ~w4198 & ~w4199;
assign w4216 = ~w4214 & w4215;
assign w4217 = ~w4196 & ~w4197;
assign w4218 = ~w4216 & w4217;
assign w4219 = ~w4194 & ~w4195;
assign w4220 = ~w4218 & w4219;
assign w4221 = ~w4193 & ~w4220;
assign w4222 = ~pi119 & pi271;
assign w4223 = pi120 & ~pi272;
assign w4224 = pi119 & ~pi271;
assign w4225 = ~pi120 & pi272;
assign w4226 = ~pi121 & pi273;
assign w4227 = pi121 & ~pi273;
assign w4228 = pi122 & ~pi274;
assign w4229 = ~pi123 & pi275;
assign w4230 = ~pi122 & pi274;
assign w4231 = pi125 & ~pi277;
assign w4232 = ~pi125 & pi277;
assign w4233 = pi126 & ~pi278;
assign w4234 = ~w4232 & w4233;
assign w4235 = ~w4231 & ~w4234;
assign w4236 = ~pi276 & ~w4235;
assign w4237 = pi123 & ~pi275;
assign w4238 = pi276 & w4235;
assign w4239 = pi124 & ~w4238;
assign w4240 = ~w4236 & ~w4237;
assign w4241 = ~w4239 & w4240;
assign w4242 = ~w4229 & ~w4230;
assign w4243 = ~w4241 & w4242;
assign w4244 = ~w4227 & ~w4228;
assign w4245 = ~w4243 & w4244;
assign w4246 = ~w4225 & ~w4226;
assign w4247 = ~w4245 & w4246;
assign w4248 = ~w4223 & ~w4224;
assign w4249 = ~w4247 & w4248;
assign w4250 = ~w4222 & ~w4249;
assign w4251 = ~w4221 & ~w4250;
assign w4252 = ~pi119 & pi247;
assign w4253 = pi120 & ~pi248;
assign w4254 = pi119 & ~pi247;
assign w4255 = ~pi120 & pi248;
assign w4256 = ~pi121 & pi249;
assign w4257 = pi121 & ~pi249;
assign w4258 = pi122 & ~pi250;
assign w4259 = pi123 & ~pi251;
assign w4260 = pi124 & ~pi252;
assign w4261 = ~pi125 & pi253;
assign w4262 = pi125 & ~pi253;
assign w4263 = pi126 & ~pi254;
assign w4264 = ~w4262 & ~w4263;
assign w4265 = ~pi124 & pi252;
assign w4266 = ~w4261 & ~w4265;
assign w4267 = ~w4264 & w4266;
assign w4268 = ~w4259 & ~w4260;
assign w4269 = ~w4267 & w4268;
assign w4270 = ~pi122 & pi250;
assign w4271 = ~pi123 & pi251;
assign w4272 = ~w4270 & ~w4271;
assign w4273 = ~w4269 & w4272;
assign w4274 = ~w4257 & ~w4258;
assign w4275 = ~w4273 & w4274;
assign w4276 = ~w4255 & ~w4256;
assign w4277 = ~w4275 & w4276;
assign w4278 = ~w4253 & ~w4254;
assign w4279 = ~w4277 & w4278;
assign w4280 = ~w4252 & ~w4279;
assign w4281 = ~w4192 & ~w4280;
assign w4282 = w4251 & w4281;
assign w4283 = ~w4134 & ~w4163;
assign w4284 = w4282 & w4283;
assign w4285 = ~pi119 & pi127;
assign w4286 = pi119 & ~pi127;
assign w4287 = pi120 & ~pi128;
assign w4288 = ~pi121 & pi129;
assign w4289 = ~pi120 & pi128;
assign w4290 = pi121 & ~pi129;
assign w4291 = pi122 & ~pi130;
assign w4292 = ~pi122 & pi130;
assign w4293 = ~pi123 & pi131;
assign w4294 = pi125 & ~pi133;
assign w4295 = ~pi125 & pi133;
assign w4296 = pi126 & ~pi134;
assign w4297 = ~w4295 & w4296;
assign w4298 = ~w4294 & ~w4297;
assign w4299 = ~pi132 & ~w4298;
assign w4300 = pi123 & ~pi131;
assign w4301 = pi132 & w4298;
assign w4302 = pi124 & ~w4301;
assign w4303 = ~w4299 & ~w4300;
assign w4304 = ~w4302 & w4303;
assign w4305 = ~w4292 & ~w4293;
assign w4306 = ~w4304 & w4305;
assign w4307 = ~w4290 & ~w4291;
assign w4308 = ~w4306 & w4307;
assign w4309 = ~w4288 & ~w4289;
assign w4310 = ~w4308 & w4309;
assign w4311 = ~w4286 & ~w4287;
assign w4312 = ~w4310 & w4311;
assign w4313 = ~w4285 & ~w4312;
assign w4314 = ~pi119 & pi167;
assign w4315 = pi119 & ~pi167;
assign w4316 = pi120 & ~pi168;
assign w4317 = pi121 & ~pi169;
assign w4318 = pi122 & ~pi170;
assign w4319 = ~pi122 & pi170;
assign w4320 = ~pi123 & pi171;
assign w4321 = pi123 & ~pi171;
assign w4322 = pi124 & ~pi172;
assign w4323 = ~pi125 & pi173;
assign w4324 = pi125 & ~pi173;
assign w4325 = pi126 & ~pi174;
assign w4326 = ~w4324 & ~w4325;
assign w4327 = ~pi124 & pi172;
assign w4328 = ~w4323 & ~w4327;
assign w4329 = ~w4326 & w4328;
assign w4330 = ~w4321 & ~w4322;
assign w4331 = ~w4329 & w4330;
assign w4332 = ~w4319 & ~w4320;
assign w4333 = ~w4331 & w4332;
assign w4334 = ~w4317 & ~w4318;
assign w4335 = ~w4333 & w4334;
assign w4336 = ~pi120 & pi168;
assign w4337 = ~pi121 & pi169;
assign w4338 = ~w4336 & ~w4337;
assign w4339 = ~w4335 & w4338;
assign w4340 = ~w4315 & ~w4316;
assign w4341 = ~w4339 & w4340;
assign w4342 = ~w4314 & ~w4341;
assign w4343 = pi119 & ~pi191;
assign w4344 = ~pi119 & pi191;
assign w4345 = pi120 & ~pi192;
assign w4346 = ~pi121 & pi193;
assign w4347 = ~pi120 & pi192;
assign w4348 = pi121 & ~pi193;
assign w4349 = pi122 & ~pi194;
assign w4350 = ~pi122 & pi194;
assign w4351 = ~pi123 & pi195;
assign w4352 = pi125 & ~pi197;
assign w4353 = ~pi125 & pi197;
assign w4354 = pi126 & ~pi198;
assign w4355 = ~w4353 & w4354;
assign w4356 = ~w4352 & ~w4355;
assign w4357 = ~pi196 & ~w4356;
assign w4358 = pi123 & ~pi195;
assign w4359 = pi196 & w4356;
assign w4360 = pi124 & ~w4359;
assign w4361 = ~w4357 & ~w4358;
assign w4362 = ~w4360 & w4361;
assign w4363 = ~w4350 & ~w4351;
assign w4364 = ~w4362 & w4363;
assign w4365 = ~w4348 & ~w4349;
assign w4366 = ~w4364 & w4365;
assign w4367 = ~w4346 & ~w4347;
assign w4368 = ~w4366 & w4367;
assign w4369 = ~w4345 & ~w4368;
assign w4370 = ~w4344 & ~w4369;
assign w4371 = ~w4343 & ~w4370;
assign w4372 = pi119 & ~pi175;
assign w4373 = ~pi119 & pi175;
assign w4374 = pi120 & ~pi176;
assign w4375 = ~pi120 & pi176;
assign w4376 = pi121 & ~pi177;
assign w4377 = ~pi121 & pi177;
assign w4378 = pi122 & ~pi178;
assign w4379 = ~pi122 & pi178;
assign w4380 = pi123 & ~pi179;
assign w4381 = ~pi123 & pi179;
assign w4382 = ~pi124 & pi180;
assign w4383 = pi125 & ~pi181;
assign w4384 = ~pi125 & pi181;
assign w4385 = pi126 & ~pi182;
assign w4386 = ~w4384 & w4385;
assign w4387 = ~w4383 & ~w4386;
assign w4388 = ~w4382 & ~w4387;
assign w4389 = pi124 & ~pi180;
assign w4390 = ~w4388 & ~w4389;
assign w4391 = ~w4381 & ~w4390;
assign w4392 = ~w4380 & ~w4391;
assign w4393 = ~w4379 & ~w4392;
assign w4394 = ~w4378 & ~w4393;
assign w4395 = ~w4377 & ~w4394;
assign w4396 = ~w4376 & ~w4395;
assign w4397 = ~w4375 & ~w4396;
assign w4398 = ~w4374 & ~w4397;
assign w4399 = ~w4373 & ~w4398;
assign w4400 = ~w4372 & ~w4399;
assign w4401 = ~w4342 & w4371;
assign w4402 = w4400 & w4401;
assign w4403 = ~pi119 & pi239;
assign w4404 = pi120 & ~pi240;
assign w4405 = pi119 & ~pi239;
assign w4406 = ~pi120 & pi240;
assign w4407 = ~pi121 & pi241;
assign w4408 = pi121 & ~pi241;
assign w4409 = pi122 & ~pi242;
assign w4410 = ~pi122 & pi242;
assign w4411 = ~pi123 & pi243;
assign w4412 = pi123 & ~pi243;
assign w4413 = pi124 & ~pi244;
assign w4414 = ~pi125 & pi245;
assign w4415 = pi125 & ~pi245;
assign w4416 = pi126 & ~pi246;
assign w4417 = ~w4415 & ~w4416;
assign w4418 = ~pi124 & pi244;
assign w4419 = ~w4414 & ~w4418;
assign w4420 = ~w4417 & w4419;
assign w4421 = ~w4412 & ~w4413;
assign w4422 = ~w4420 & w4421;
assign w4423 = ~w4410 & ~w4411;
assign w4424 = ~w4422 & w4423;
assign w4425 = ~w4408 & ~w4409;
assign w4426 = ~w4424 & w4425;
assign w4427 = ~w4406 & ~w4407;
assign w4428 = ~w4426 & w4427;
assign w4429 = ~w4404 & ~w4405;
assign w4430 = ~w4428 & w4429;
assign w4431 = ~w4403 & ~w4430;
assign w4432 = ~pi119 & pi231;
assign w4433 = ~pi121 & pi233;
assign w4434 = ~pi120 & pi232;
assign w4435 = pi121 & ~pi233;
assign w4436 = pi122 & ~pi234;
assign w4437 = ~pi122 & pi234;
assign w4438 = ~pi123 & pi235;
assign w4439 = pi125 & ~pi237;
assign w4440 = ~pi125 & pi237;
assign w4441 = pi126 & ~pi238;
assign w4442 = ~w4440 & w4441;
assign w4443 = ~w4439 & ~w4442;
assign w4444 = ~pi236 & ~w4443;
assign w4445 = pi123 & ~pi235;
assign w4446 = pi236 & w4443;
assign w4447 = pi124 & ~w4446;
assign w4448 = ~w4444 & ~w4445;
assign w4449 = ~w4447 & w4448;
assign w4450 = ~w4437 & ~w4438;
assign w4451 = ~w4449 & w4450;
assign w4452 = ~w4435 & ~w4436;
assign w4453 = ~w4451 & w4452;
assign w4454 = ~w4433 & ~w4434;
assign w4455 = ~w4453 & w4454;
assign w4456 = pi119 & ~pi231;
assign w4457 = pi120 & ~pi232;
assign w4458 = ~w4456 & ~w4457;
assign w4459 = ~w4455 & w4458;
assign w4460 = ~w4432 & ~w4459;
assign w4461 = ~w4431 & ~w4460;
assign w4462 = ~pi119 & pi151;
assign w4463 = pi120 & ~pi152;
assign w4464 = pi119 & ~pi151;
assign w4465 = ~pi120 & pi152;
assign w4466 = ~pi121 & pi153;
assign w4467 = pi121 & ~pi153;
assign w4468 = pi122 & ~pi154;
assign w4469 = pi123 & ~pi155;
assign w4470 = pi124 & ~pi156;
assign w4471 = ~pi125 & pi157;
assign w4472 = pi125 & ~pi157;
assign w4473 = pi126 & ~pi158;
assign w4474 = ~w4472 & ~w4473;
assign w4475 = ~pi124 & pi156;
assign w4476 = ~w4471 & ~w4475;
assign w4477 = ~w4474 & w4476;
assign w4478 = ~w4469 & ~w4470;
assign w4479 = ~w4477 & w4478;
assign w4480 = ~pi122 & pi154;
assign w4481 = ~pi123 & pi155;
assign w4482 = ~w4480 & ~w4481;
assign w4483 = ~w4479 & w4482;
assign w4484 = ~w4467 & ~w4468;
assign w4485 = ~w4483 & w4484;
assign w4486 = ~w4465 & ~w4466;
assign w4487 = ~w4485 & w4486;
assign w4488 = ~w4463 & ~w4464;
assign w4489 = ~w4487 & w4488;
assign w4490 = ~w4462 & ~w4489;
assign w4491 = pi119 & ~pi159;
assign w4492 = ~pi119 & pi159;
assign w4493 = pi120 & ~pi160;
assign w4494 = ~pi120 & pi160;
assign w4495 = pi121 & ~pi161;
assign w4496 = ~pi121 & pi161;
assign w4497 = pi122 & ~pi162;
assign w4498 = ~pi122 & pi162;
assign w4499 = pi123 & ~pi163;
assign w4500 = ~pi123 & pi163;
assign w4501 = ~pi124 & pi164;
assign w4502 = pi125 & ~pi165;
assign w4503 = ~pi125 & pi165;
assign w4504 = pi126 & ~pi166;
assign w4505 = ~w4503 & w4504;
assign w4506 = ~w4502 & ~w4505;
assign w4507 = ~w4501 & ~w4506;
assign w4508 = pi124 & ~pi164;
assign w4509 = ~w4507 & ~w4508;
assign w4510 = ~w4500 & ~w4509;
assign w4511 = ~w4499 & ~w4510;
assign w4512 = ~w4498 & ~w4511;
assign w4513 = ~w4497 & ~w4512;
assign w4514 = ~w4496 & ~w4513;
assign w4515 = ~w4495 & ~w4514;
assign w4516 = ~w4494 & ~w4515;
assign w4517 = ~w4493 & ~w4516;
assign w4518 = ~w4492 & ~w4517;
assign w4519 = ~w4491 & ~w4518;
assign w4520 = w4461 & ~w4490;
assign w4521 = w4519 & w4520;
assign w4522 = w4402 & w4521;
assign w4523 = ~pi119 & pi183;
assign w4524 = pi119 & ~pi183;
assign w4525 = pi120 & ~pi184;
assign w4526 = ~pi120 & pi184;
assign w4527 = ~pi121 & pi185;
assign w4528 = pi121 & ~pi185;
assign w4529 = pi122 & ~pi186;
assign w4530 = pi123 & ~pi187;
assign w4531 = pi124 & ~pi188;
assign w4532 = ~pi125 & pi189;
assign w4533 = pi125 & ~pi189;
assign w4534 = pi126 & ~pi190;
assign w4535 = ~w4533 & ~w4534;
assign w4536 = ~pi124 & pi188;
assign w4537 = ~w4532 & ~w4536;
assign w4538 = ~w4535 & w4537;
assign w4539 = ~w4530 & ~w4531;
assign w4540 = ~w4538 & w4539;
assign w4541 = ~pi122 & pi186;
assign w4542 = ~pi123 & pi187;
assign w4543 = ~w4541 & ~w4542;
assign w4544 = ~w4540 & w4543;
assign w4545 = ~w4528 & ~w4529;
assign w4546 = ~w4544 & w4545;
assign w4547 = ~w4526 & ~w4527;
assign w4548 = ~w4546 & w4547;
assign w4549 = ~w4524 & ~w4525;
assign w4550 = ~w4548 & w4549;
assign w4551 = ~w4523 & ~w4550;
assign w4552 = ~pi119 & pi223;
assign w4553 = pi120 & ~pi224;
assign w4554 = pi119 & ~pi223;
assign w4555 = ~pi120 & pi224;
assign w4556 = ~pi121 & pi225;
assign w4557 = pi121 & ~pi225;
assign w4558 = pi122 & ~pi226;
assign w4559 = pi123 & ~pi227;
assign w4560 = pi124 & ~pi228;
assign w4561 = ~pi125 & pi229;
assign w4562 = pi125 & ~pi229;
assign w4563 = pi126 & ~pi230;
assign w4564 = ~w4562 & ~w4563;
assign w4565 = ~pi124 & pi228;
assign w4566 = ~w4561 & ~w4565;
assign w4567 = ~w4564 & w4566;
assign w4568 = ~w4559 & ~w4560;
assign w4569 = ~w4567 & w4568;
assign w4570 = ~pi122 & pi226;
assign w4571 = ~pi123 & pi227;
assign w4572 = ~w4570 & ~w4571;
assign w4573 = ~w4569 & w4572;
assign w4574 = ~w4557 & ~w4558;
assign w4575 = ~w4573 & w4574;
assign w4576 = ~w4555 & ~w4556;
assign w4577 = ~w4575 & w4576;
assign w4578 = ~w4553 & ~w4554;
assign w4579 = ~w4577 & w4578;
assign w4580 = ~w4552 & ~w4579;
assign w4581 = ~pi119 & pi207;
assign w4582 = pi119 & ~pi207;
assign w4583 = pi120 & ~pi208;
assign w4584 = ~pi120 & pi208;
assign w4585 = ~pi121 & pi209;
assign w4586 = pi121 & ~pi209;
assign w4587 = pi122 & ~pi210;
assign w4588 = ~pi122 & pi210;
assign w4589 = ~pi123 & pi211;
assign w4590 = pi123 & ~pi211;
assign w4591 = pi124 & ~pi212;
assign w4592 = ~pi125 & pi213;
assign w4593 = pi125 & ~pi213;
assign w4594 = pi126 & ~pi214;
assign w4595 = ~w4593 & ~w4594;
assign w4596 = ~pi124 & pi212;
assign w4597 = ~w4592 & ~w4596;
assign w4598 = ~w4595 & w4597;
assign w4599 = ~w4590 & ~w4591;
assign w4600 = ~w4598 & w4599;
assign w4601 = ~w4588 & ~w4589;
assign w4602 = ~w4600 & w4601;
assign w4603 = ~w4586 & ~w4587;
assign w4604 = ~w4602 & w4603;
assign w4605 = ~w4584 & ~w4585;
assign w4606 = ~w4604 & w4605;
assign w4607 = ~w4582 & ~w4583;
assign w4608 = ~w4606 & w4607;
assign w4609 = ~w4581 & ~w4608;
assign w4610 = ~pi119 & pi199;
assign w4611 = pi120 & ~pi200;
assign w4612 = pi119 & ~pi199;
assign w4613 = pi121 & ~pi201;
assign w4614 = pi122 & ~pi202;
assign w4615 = ~pi122 & pi202;
assign w4616 = ~pi123 & pi203;
assign w4617 = pi123 & ~pi203;
assign w4618 = pi124 & ~pi204;
assign w4619 = ~pi125 & pi205;
assign w4620 = pi125 & ~pi205;
assign w4621 = pi126 & ~pi206;
assign w4622 = ~w4620 & ~w4621;
assign w4623 = ~pi124 & pi204;
assign w4624 = ~w4619 & ~w4623;
assign w4625 = ~w4622 & w4624;
assign w4626 = ~w4617 & ~w4618;
assign w4627 = ~w4625 & w4626;
assign w4628 = ~w4615 & ~w4616;
assign w4629 = ~w4627 & w4628;
assign w4630 = ~w4613 & ~w4614;
assign w4631 = ~w4629 & w4630;
assign w4632 = ~pi120 & pi200;
assign w4633 = ~pi121 & pi201;
assign w4634 = ~w4632 & ~w4633;
assign w4635 = ~w4631 & w4634;
assign w4636 = ~w4611 & ~w4612;
assign w4637 = ~w4635 & w4636;
assign w4638 = ~w4610 & ~w4637;
assign w4639 = ~pi119 & pi215;
assign w4640 = pi120 & ~pi216;
assign w4641 = pi119 & ~pi215;
assign w4642 = ~pi120 & pi216;
assign w4643 = ~pi121 & pi217;
assign w4644 = pi121 & ~pi217;
assign w4645 = pi122 & ~pi218;
assign w4646 = pi123 & ~pi219;
assign w4647 = pi124 & ~pi220;
assign w4648 = ~pi125 & pi221;
assign w4649 = pi125 & ~pi221;
assign w4650 = pi126 & ~pi222;
assign w4651 = ~w4649 & ~w4650;
assign w4652 = ~pi124 & pi220;
assign w4653 = ~w4648 & ~w4652;
assign w4654 = ~w4651 & w4653;
assign w4655 = ~w4646 & ~w4647;
assign w4656 = ~w4654 & w4655;
assign w4657 = ~pi122 & pi218;
assign w4658 = ~pi123 & pi219;
assign w4659 = ~w4657 & ~w4658;
assign w4660 = ~w4656 & w4659;
assign w4661 = ~w4644 & ~w4645;
assign w4662 = ~w4660 & w4661;
assign w4663 = ~w4642 & ~w4643;
assign w4664 = ~w4662 & w4663;
assign w4665 = ~w4640 & ~w4641;
assign w4666 = ~w4664 & w4665;
assign w4667 = ~w4639 & ~w4666;
assign w4668 = ~w4609 & ~w4638;
assign w4669 = ~w4667 & w4668;
assign w4670 = ~w4580 & w4669;
assign w4671 = ~w4551 & w4670;
assign w4672 = w4522 & w4671;
assign w4673 = w2753 & ~w3296;
assign w4674 = (w4673 & ~w3399) | (w4673 & w17009) | (~w3399 & w17009);
assign w4675 = w754 & w3350;
assign w4676 = (w4675 & ~w3419) | (w4675 & w17010) | (~w3419 & w17010);
assign w4677 = ~w2540 & ~w3306;
assign w4678 = ~w2473 & w4677;
assign w4679 = ~w3387 & w4678;
assign w4680 = w4071 & ~w4313;
assign w4681 = w4284 & w4680;
assign w4682 = w4672 & w4681;
assign w4683 = ~w4105 & w4682;
assign w4684 = ~w4674 & w4683;
assign w4685 = ~w4676 & ~w4679;
assign w4686 = w4684 & w4685;
assign w4687 = w4685 & w18320;
assign w4688 = pi011 & w4687;
assign w4689 = w3392 & ~w4094;
assign w4690 = ~w3387 & w3394;
assign w4691 = (~w2632 & ~w4082) | (~w2632 & w17011) | (~w4082 & w17011);
assign w4692 = w3258 & w4691;
assign w4693 = ~w4689 & ~w4690;
assign w4694 = ~w4692 & w4693;
assign w4695 = ~w2667 & ~w4051;
assign w4696 = (w3389 & ~w3419) | (w3389 & w17012) | (~w3419 & w17012);
assign w4697 = ~w4695 & ~w4696;
assign w4698 = w3287 & ~w4071;
assign w4699 = w2754 & ~w4698;
assign w4700 = w3390 & w4699;
assign w4701 = w3349 & w16247;
assign w4702 = ~w3402 & w4701;
assign w4703 = w3257 & w4702;
assign w4704 = w4697 & w4703;
assign w4705 = w4694 & w4704;
assign w4706 = pi007 & w4705;
assign w4707 = ~w3977 & ~w4036;
assign w4708 = w2542 & w4060;
assign w4709 = ~w1249 & w1253;
assign w4710 = ~w1245 & w4709;
assign w4711 = w1259 & ~w4710;
assign w4712 = w310 & ~w4711;
assign w4713 = w4708 & w4712;
assign w4714 = pi103 & pi119;
assign w4715 = pi127 & ~w4714;
assign w4716 = ~w851 & ~w4054;
assign w4717 = ~w2532 & w4716;
assign w4718 = w2218 & w2222;
assign w4719 = w2227 & ~w4718;
assign w4720 = ~w2988 & ~w4719;
assign w4721 = w2627 & w4720;
assign w4722 = w4717 & w4721;
assign w4723 = ~w344 & ~w693;
assign w4724 = pi071 & pi087;
assign w4725 = pi127 & ~w4724;
assign w4726 = ~w823 & ~w4725;
assign w4727 = ~w1170 & w4723;
assign w4728 = w4726 & w4727;
assign w4729 = w436 & ~w2545;
assign w4730 = ~w1250 & ~w1360;
assign w4731 = ~w407 & w4730;
assign w4732 = ~w951 & w4731;
assign w4733 = w4057 & w4732;
assign w4734 = w4728 & w4733;
assign w4735 = w4729 & w4734;
assign w4736 = w29 & ~w4715;
assign w4737 = w4735 & w4736;
assign w4738 = w4713 & w4737;
assign w4739 = w4722 & w4738;
assign w4740 = w4062 & w4707;
assign w4741 = w4739 & w4740;
assign w4742 = ~w4312 & w4741;
assign w4743 = pi012 & w4742;
assign w4744 = (w4043 & ~w3419) | (w4043 & w17013) | (~w3419 & w17013);
assign w4745 = w4038 & ~w4071;
assign w4746 = w3745 & ~w4745;
assign w4747 = w4105 & w4746;
assign w4748 = ~w4744 & w4747;
assign w4749 = w2667 & ~w3296;
assign w4750 = (w4749 & ~w3399) | (w4749 & w17014) | (~w3399 & w17014);
assign w4751 = w4041 & ~w4094;
assign w4752 = ~w3387 & w4040;
assign w4753 = ~w4691 & ~w4750;
assign w4754 = ~w4751 & ~w4752;
assign w4755 = w4753 & w4754;
assign w4756 = w3980 & w4748;
assign w4757 = w4755 & w4756;
assign w4758 = pi009 & w4757;
assign w4759 = (w4075 & ~w3419) | (w4075 & w17549) | (~w3419 & w17549);
assign w4760 = (w4076 & ~w3399) | (w4076 & w17550) | (~w3399 & w17550);
assign w4761 = ~w3387 & w4078;
assign w4762 = w4073 & ~w4094;
assign w4763 = w3352 & ~w4760;
assign w4764 = ~w4761 & ~w4762;
assign w4765 = w4763 & w4764;
assign w4766 = w4691 & ~w4759;
assign w4767 = w4765 & w4766;
assign w4768 = pi008 & w4767;
assign w4769 = ~w3387 & w4677;
assign w4770 = ~w3387 & w17015;
assign w4771 = (~w4038 & ~w4050) | (~w4038 & w17016) | (~w4050 & w17016);
assign w4772 = w1388 & w3391;
assign w4773 = ~w4094 & w4772;
assign w4774 = (~w3296 & ~w3399) | (~w3296 & w17017) | (~w3399 & w17017);
assign w4775 = ~w3287 & w4774;
assign w4776 = w723 & w3350;
assign w4777 = (w4776 & ~w3419) | (w4776 & w17018) | (~w3419 & w17018);
assign w4778 = ~w4071 & ~w4771;
assign w4779 = ~w4691 & w4778;
assign w4780 = ~w4773 & ~w4777;
assign w4781 = w4779 & w4780;
assign w4782 = ~w4770 & ~w4775;
assign w4783 = w4781 & w4782;
assign w4784 = pi010 & w4783;
assign w4785 = ~pi005 & ~w1949;
assign w4786 = w3377 & ~w4094;
assign w4787 = (w3372 & ~w3399) | (w3372 & w17019) | (~w3399 & w17019);
assign w4788 = (w3380 & ~w4082) | (w3380 & w17020) | (~w4082 & w17020);
assign w4789 = (w3373 & ~w3419) | (w3373 & w17021) | (~w3419 & w17021);
assign w4790 = ~w4786 & ~w4787;
assign w4791 = ~w4788 & ~w4789;
assign w4792 = w4790 & w4791;
assign w4793 = (w2502 & ~w4050) | (w2502 & w17022) | (~w4050 & w17022);
assign w4794 = w2260 & ~w4071;
assign w4795 = w2322 & w2445;
assign w4796 = ~w2291 & w4795;
assign w4797 = (w3371 & ~w3349) | (w3371 & w16248) | (~w3349 & w16248);
assign w4798 = w2230 & ~w2473;
assign w4799 = w4796 & w4798;
assign w4800 = ~w4794 & w4799;
assign w4801 = w3379 & w4800;
assign w4802 = w3376 & w4801;
assign w4803 = ~w3387 & w4802;
assign w4804 = ~w4793 & ~w4797;
assign w4805 = w4803 & w4804;
assign w4806 = w4792 & w4805;
assign w4807 = w4785 & w4806;
assign w4808 = (w3361 & ~w3349) | (w3361 & w16249) | (~w3349 & w16249);
assign w4809 = w3362 & ~w4808;
assign w4810 = w4102 & w4809;
assign w4811 = w3360 & ~w4082;
assign w4812 = (w1417 & ~w4050) | (w1417 & w17023) | (~w4050 & w17023);
assign w4813 = w3359 & ~w3387;
assign w4814 = ~w1388 & ~w4071;
assign w4815 = w1169 & w1670;
assign w4816 = w3314 & w4815;
assign w4817 = w1293 & w1756;
assign w4818 = w4816 & w4817;
assign w4819 = ~w4814 & w4818;
assign w4820 = ~w3356 & w4819;
assign w4821 = w3405 & w4819;
assign w4822 = (~w4820 & ~w3419) | (~w4820 & w17024) | (~w3419 & w17024);
assign w4823 = (w3357 & ~w3399) | (w3357 & w17551) | (~w3399 & w17551);
assign w4824 = ~w4811 & ~w4812;
assign w4825 = ~w4813 & w4824;
assign w4826 = ~w4822 & ~w4823;
assign w4827 = w4825 & w4826;
assign w4828 = w4810 & w4827;
assign w4829 = pi003 & w4828;
assign w4830 = w4803 & w17025;
assign w4831 = w4792 & w4830;
assign w4832 = ~w3387 & w3406;
assign w4833 = (w278 & ~w4050) | (w278 & w17026) | (~w4050 & w17026);
assign w4834 = ~w723 & ~w4070;
assign w4835 = w220 & w597;
assign w4836 = w249 & w692;
assign w4837 = w4835 & w4836;
assign w4838 = w914 & w4837;
assign w4839 = w822 & w4838;
assign w4840 = w754 & w4839;
assign w4841 = ~w4834 & w4840;
assign w4842 = ~w4833 & w4841;
assign w4843 = ~w4832 & w4842;
assign w4844 = (w3409 & ~w4082) | (w3409 & w17027) | (~w4082 & w17027);
assign w4845 = (w3408 & ~w3399) | (w3408 & w17028) | (~w3399 & w17028);
assign w4846 = w3407 & ~w4094;
assign w4847 = (~w373 & ~w3348) | (~w373 & w16250) | (~w3348 & w16250);
assign w4848 = w2634 & ~w4847;
assign w4849 = ~w3420 & w4848;
assign w4850 = ~w4844 & ~w4845;
assign w4851 = ~w4846 & w4849;
assign w4852 = w4850 & w4851;
assign w4853 = ~w4832 & w17029;
assign w4854 = w4852 & w4853;
assign w4855 = pi001 & w4854;
assign w4856 = ~w4829 & ~w4831;
assign w4857 = ~w4855 & w4856;
assign w4858 = ~w4100 & ~w4807;
assign w4859 = ~w4857 & w4858;
assign w4860 = ~w4101 & ~w4743;
assign w4861 = ~w4688 & w4860;
assign w4862 = ~w4706 & ~w4758;
assign w4863 = ~w4768 & ~w4784;
assign w4864 = w4862 & w4863;
assign w4865 = w4861 & w4864;
assign w4866 = ~w4859 & w4865;
assign w4867 = ~pi135 & pi207;
assign w4868 = pi136 & ~pi208;
assign w4869 = pi135 & ~pi207;
assign w4870 = ~pi136 & pi208;
assign w4871 = ~pi137 & pi209;
assign w4872 = pi137 & ~pi209;
assign w4873 = pi138 & ~pi210;
assign w4874 = ~pi138 & pi210;
assign w4875 = ~pi139 & pi211;
assign w4876 = pi139 & ~pi211;
assign w4877 = pi140 & ~pi212;
assign w4878 = ~pi141 & pi213;
assign w4879 = pi141 & ~pi213;
assign w4880 = pi142 & ~pi214;
assign w4881 = ~w4879 & ~w4880;
assign w4882 = ~pi140 & pi212;
assign w4883 = ~w4878 & ~w4882;
assign w4884 = ~w4881 & w4883;
assign w4885 = ~w4876 & ~w4877;
assign w4886 = ~w4884 & w4885;
assign w4887 = ~w4874 & ~w4875;
assign w4888 = ~w4886 & w4887;
assign w4889 = ~w4872 & ~w4873;
assign w4890 = ~w4888 & w4889;
assign w4891 = ~w4870 & ~w4871;
assign w4892 = ~w4890 & w4891;
assign w4893 = ~w4868 & ~w4869;
assign w4894 = ~w4892 & w4893;
assign w4895 = ~w4867 & ~w4894;
assign w4896 = ~pi135 & pi199;
assign w4897 = pi135 & ~pi199;
assign w4898 = pi136 & ~pi200;
assign w4899 = ~pi136 & pi200;
assign w4900 = ~pi137 & pi201;
assign w4901 = pi137 & ~pi201;
assign w4902 = pi138 & ~pi202;
assign w4903 = pi139 & ~pi203;
assign w4904 = pi140 & ~pi204;
assign w4905 = ~pi141 & pi205;
assign w4906 = pi141 & ~pi205;
assign w4907 = pi142 & ~pi206;
assign w4908 = ~w4906 & ~w4907;
assign w4909 = ~pi140 & pi204;
assign w4910 = ~w4905 & ~w4909;
assign w4911 = ~w4908 & w4910;
assign w4912 = ~w4903 & ~w4904;
assign w4913 = ~w4911 & w4912;
assign w4914 = ~pi138 & pi202;
assign w4915 = ~pi139 & pi203;
assign w4916 = ~w4914 & ~w4915;
assign w4917 = ~w4913 & w4916;
assign w4918 = ~w4901 & ~w4902;
assign w4919 = ~w4917 & w4918;
assign w4920 = ~w4899 & ~w4900;
assign w4921 = ~w4919 & w4920;
assign w4922 = ~w4897 & ~w4898;
assign w4923 = ~w4921 & w4922;
assign w4924 = ~w4896 & ~w4923;
assign w4925 = ~w4895 & ~w4924;
assign w4926 = ~pi135 & pi271;
assign w4927 = pi136 & ~pi272;
assign w4928 = pi135 & ~pi271;
assign w4929 = pi137 & ~pi273;
assign w4930 = pi138 & ~pi274;
assign w4931 = ~pi138 & pi274;
assign w4932 = ~pi139 & pi275;
assign w4933 = pi139 & ~pi275;
assign w4934 = pi140 & ~pi276;
assign w4935 = ~pi141 & pi277;
assign w4936 = pi141 & ~pi277;
assign w4937 = pi142 & ~pi278;
assign w4938 = ~w4936 & ~w4937;
assign w4939 = ~pi140 & pi276;
assign w4940 = ~w4935 & ~w4939;
assign w4941 = ~w4938 & w4940;
assign w4942 = ~w4933 & ~w4934;
assign w4943 = ~w4941 & w4942;
assign w4944 = ~w4931 & ~w4932;
assign w4945 = ~w4943 & w4944;
assign w4946 = ~w4929 & ~w4930;
assign w4947 = ~w4945 & w4946;
assign w4948 = ~pi136 & pi272;
assign w4949 = ~pi137 & pi273;
assign w4950 = ~w4948 & ~w4949;
assign w4951 = ~w4947 & w4950;
assign w4952 = ~w4927 & ~w4928;
assign w4953 = ~w4951 & w4952;
assign w4954 = ~w4926 & ~w4953;
assign w4955 = ~pi135 & pi263;
assign w4956 = pi135 & ~pi263;
assign w4957 = pi136 & ~pi264;
assign w4958 = ~pi136 & pi264;
assign w4959 = ~pi137 & pi265;
assign w4960 = pi137 & ~pi265;
assign w4961 = pi138 & ~pi266;
assign w4962 = pi139 & ~pi267;
assign w4963 = pi140 & ~pi268;
assign w4964 = ~pi141 & pi269;
assign w4965 = pi141 & ~pi269;
assign w4966 = pi142 & ~pi270;
assign w4967 = ~w4965 & ~w4966;
assign w4968 = ~pi140 & pi268;
assign w4969 = ~w4964 & ~w4968;
assign w4970 = ~w4967 & w4969;
assign w4971 = ~w4962 & ~w4963;
assign w4972 = ~w4970 & w4971;
assign w4973 = ~pi138 & pi266;
assign w4974 = ~pi139 & pi267;
assign w4975 = ~w4973 & ~w4974;
assign w4976 = ~w4972 & w4975;
assign w4977 = ~w4960 & ~w4961;
assign w4978 = ~w4976 & w4977;
assign w4979 = ~w4958 & ~w4959;
assign w4980 = ~w4978 & w4979;
assign w4981 = ~w4956 & ~w4957;
assign w4982 = ~w4980 & w4981;
assign w4983 = ~w4955 & ~w4982;
assign w4984 = ~w4954 & ~w4983;
assign w4985 = ~pi135 & pi215;
assign w4986 = pi136 & ~pi216;
assign w4987 = pi135 & ~pi215;
assign w4988 = ~pi136 & pi216;
assign w4989 = ~pi137 & pi217;
assign w4990 = pi137 & ~pi217;
assign w4991 = pi138 & ~pi218;
assign w4992 = ~pi138 & pi218;
assign w4993 = ~pi139 & pi219;
assign w4994 = pi139 & ~pi219;
assign w4995 = pi140 & ~pi220;
assign w4996 = ~pi141 & pi221;
assign w4997 = pi141 & ~pi221;
assign w4998 = pi142 & ~pi222;
assign w4999 = ~w4997 & ~w4998;
assign w5000 = ~pi140 & pi220;
assign w5001 = ~w4996 & ~w5000;
assign w5002 = ~w4999 & w5001;
assign w5003 = ~w4994 & ~w4995;
assign w5004 = ~w5002 & w5003;
assign w5005 = ~w4992 & ~w4993;
assign w5006 = ~w5004 & w5005;
assign w5007 = ~w4990 & ~w4991;
assign w5008 = ~w5006 & w5007;
assign w5009 = ~w4988 & ~w4989;
assign w5010 = ~w5008 & w5009;
assign w5011 = ~w4986 & ~w4987;
assign w5012 = ~w5010 & w5011;
assign w5013 = ~w4985 & ~w5012;
assign w5014 = ~pi135 & pi223;
assign w5015 = pi135 & ~pi223;
assign w5016 = pi136 & ~pi224;
assign w5017 = pi137 & ~pi225;
assign w5018 = pi138 & ~pi226;
assign w5019 = ~pi138 & pi226;
assign w5020 = ~pi139 & pi227;
assign w5021 = pi139 & ~pi227;
assign w5022 = pi140 & ~pi228;
assign w5023 = ~pi141 & pi229;
assign w5024 = pi141 & ~pi229;
assign w5025 = pi142 & ~pi230;
assign w5026 = ~w5024 & ~w5025;
assign w5027 = ~pi140 & pi228;
assign w5028 = ~w5023 & ~w5027;
assign w5029 = ~w5026 & w5028;
assign w5030 = ~w5021 & ~w5022;
assign w5031 = ~w5029 & w5030;
assign w5032 = ~w5019 & ~w5020;
assign w5033 = ~w5031 & w5032;
assign w5034 = ~w5017 & ~w5018;
assign w5035 = ~w5033 & w5034;
assign w5036 = ~pi136 & pi224;
assign w5037 = ~pi137 & pi225;
assign w5038 = ~w5036 & ~w5037;
assign w5039 = ~w5035 & w5038;
assign w5040 = ~w5015 & ~w5016;
assign w5041 = ~w5039 & w5040;
assign w5042 = ~w5014 & ~w5041;
assign w5043 = ~pi135 & pi255;
assign w5044 = pi136 & ~pi256;
assign w5045 = pi135 & ~pi255;
assign w5046 = ~pi136 & pi256;
assign w5047 = ~pi137 & pi257;
assign w5048 = pi137 & ~pi257;
assign w5049 = pi138 & ~pi258;
assign w5050 = ~pi139 & pi259;
assign w5051 = ~pi138 & pi258;
assign w5052 = pi141 & ~pi261;
assign w5053 = ~pi141 & pi261;
assign w5054 = pi142 & ~pi262;
assign w5055 = ~w5053 & w5054;
assign w5056 = ~w5052 & ~w5055;
assign w5057 = ~pi260 & ~w5056;
assign w5058 = pi139 & ~pi259;
assign w5059 = pi260 & w5056;
assign w5060 = pi140 & ~w5059;
assign w5061 = ~w5057 & ~w5058;
assign w5062 = ~w5060 & w5061;
assign w5063 = ~w5050 & ~w5051;
assign w5064 = ~w5062 & w5063;
assign w5065 = ~w5048 & ~w5049;
assign w5066 = ~w5064 & w5065;
assign w5067 = ~w5046 & ~w5047;
assign w5068 = ~w5066 & w5067;
assign w5069 = ~w5044 & ~w5045;
assign w5070 = ~w5068 & w5069;
assign w5071 = ~w5043 & ~w5070;
assign w5072 = ~pi135 & pi231;
assign w5073 = pi135 & ~pi231;
assign w5074 = pi136 & ~pi232;
assign w5075 = ~pi136 & pi232;
assign w5076 = ~pi137 & pi233;
assign w5077 = pi137 & ~pi233;
assign w5078 = pi138 & ~pi234;
assign w5079 = pi139 & ~pi235;
assign w5080 = pi140 & ~pi236;
assign w5081 = ~pi141 & pi237;
assign w5082 = pi141 & ~pi237;
assign w5083 = pi142 & ~pi238;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = ~pi140 & pi236;
assign w5086 = ~w5081 & ~w5085;
assign w5087 = ~w5084 & w5086;
assign w5088 = ~w5079 & ~w5080;
assign w5089 = ~w5087 & w5088;
assign w5090 = ~pi138 & pi234;
assign w5091 = ~pi139 & pi235;
assign w5092 = ~w5090 & ~w5091;
assign w5093 = ~w5089 & w5092;
assign w5094 = ~w5077 & ~w5078;
assign w5095 = ~w5093 & w5094;
assign w5096 = ~w5075 & ~w5076;
assign w5097 = ~w5095 & w5096;
assign w5098 = ~w5073 & ~w5074;
assign w5099 = ~w5097 & w5098;
assign w5100 = ~w5072 & ~w5099;
assign w5101 = ~pi135 & pi239;
assign w5102 = pi136 & ~pi240;
assign w5103 = pi135 & ~pi239;
assign w5104 = ~pi136 & pi240;
assign w5105 = ~pi137 & pi241;
assign w5106 = pi137 & ~pi241;
assign w5107 = pi138 & ~pi242;
assign w5108 = ~pi138 & pi242;
assign w5109 = ~pi139 & pi243;
assign w5110 = pi139 & ~pi243;
assign w5111 = pi140 & ~pi244;
assign w5112 = ~pi141 & pi245;
assign w5113 = pi141 & ~pi245;
assign w5114 = pi142 & ~pi246;
assign w5115 = ~w5113 & ~w5114;
assign w5116 = ~pi140 & pi244;
assign w5117 = ~w5112 & ~w5116;
assign w5118 = ~w5115 & w5117;
assign w5119 = ~w5110 & ~w5111;
assign w5120 = ~w5118 & w5119;
assign w5121 = ~w5108 & ~w5109;
assign w5122 = ~w5120 & w5121;
assign w5123 = ~w5106 & ~w5107;
assign w5124 = ~w5122 & w5123;
assign w5125 = ~w5104 & ~w5105;
assign w5126 = ~w5124 & w5125;
assign w5127 = ~w5102 & ~w5103;
assign w5128 = ~w5126 & w5127;
assign w5129 = ~w5101 & ~w5128;
assign w5130 = ~pi135 & pi247;
assign w5131 = pi135 & ~pi247;
assign w5132 = ~pi136 & pi248;
assign w5133 = pi136 & ~pi248;
assign w5134 = ~pi137 & pi249;
assign w5135 = pi137 & ~pi249;
assign w5136 = pi138 & ~pi250;
assign w5137 = ~pi138 & pi250;
assign w5138 = ~pi139 & pi251;
assign w5139 = pi141 & ~pi253;
assign w5140 = ~pi141 & pi253;
assign w5141 = pi142 & ~pi254;
assign w5142 = ~w5140 & w5141;
assign w5143 = ~w5139 & ~w5142;
assign w5144 = ~pi252 & ~w5143;
assign w5145 = pi139 & ~pi251;
assign w5146 = pi252 & w5143;
assign w5147 = pi140 & ~w5146;
assign w5148 = ~w5144 & ~w5145;
assign w5149 = ~w5147 & w5148;
assign w5150 = ~w5137 & ~w5138;
assign w5151 = ~w5149 & w5150;
assign w5152 = ~w5135 & ~w5136;
assign w5153 = ~w5151 & w5152;
assign w5154 = ~w5134 & ~w5153;
assign w5155 = ~w5133 & ~w5154;
assign w5156 = ~w5132 & ~w5155;
assign w5157 = ~w5131 & ~w5156;
assign w5158 = ~w5130 & ~w5157;
assign w5159 = ~w5100 & ~w5129;
assign w5160 = ~w5071 & w5159;
assign w5161 = ~w5158 & w5160;
assign w5162 = ~w5042 & w5161;
assign w5163 = ~w5013 & w5162;
assign w5164 = pi135 & ~pi183;
assign w5165 = ~pi135 & pi183;
assign w5166 = pi136 & ~pi184;
assign w5167 = ~pi136 & pi184;
assign w5168 = pi137 & ~pi185;
assign w5169 = ~pi137 & pi185;
assign w5170 = pi138 & ~pi186;
assign w5171 = ~pi138 & pi186;
assign w5172 = pi139 & ~pi187;
assign w5173 = ~pi139 & pi187;
assign w5174 = ~pi140 & pi188;
assign w5175 = pi141 & ~pi189;
assign w5176 = ~pi141 & pi189;
assign w5177 = pi142 & ~pi190;
assign w5178 = ~w5176 & w5177;
assign w5179 = ~w5175 & ~w5178;
assign w5180 = ~w5174 & ~w5179;
assign w5181 = pi140 & ~pi188;
assign w5182 = ~w5180 & ~w5181;
assign w5183 = ~w5173 & ~w5182;
assign w5184 = ~w5172 & ~w5183;
assign w5185 = ~w5171 & ~w5184;
assign w5186 = ~w5170 & ~w5185;
assign w5187 = ~w5169 & ~w5186;
assign w5188 = ~w5168 & ~w5187;
assign w5189 = ~w5167 & ~w5188;
assign w5190 = ~w5166 & ~w5189;
assign w5191 = ~w5165 & ~w5190;
assign w5192 = ~w5164 & ~w5191;
assign w5193 = w4925 & w4984;
assign w5194 = w5192 & w5193;
assign w5195 = w5163 & w5194;
assign w5196 = ~pi135 & pi159;
assign w5197 = pi135 & ~pi159;
assign w5198 = ~pi136 & pi160;
assign w5199 = pi136 & ~pi160;
assign w5200 = ~pi137 & pi161;
assign w5201 = pi137 & ~pi161;
assign w5202 = pi138 & ~pi162;
assign w5203 = ~pi139 & pi163;
assign w5204 = ~pi138 & pi162;
assign w5205 = pi139 & ~pi163;
assign w5206 = pi140 & ~pi164;
assign w5207 = ~pi140 & pi164;
assign w5208 = pi141 & ~pi165;
assign w5209 = ~pi141 & pi165;
assign w5210 = pi142 & ~pi166;
assign w5211 = ~w5209 & w5210;
assign w5212 = ~w5208 & ~w5211;
assign w5213 = ~w5207 & ~w5212;
assign w5214 = ~w5205 & ~w5206;
assign w5215 = ~w5213 & w5214;
assign w5216 = ~w5203 & ~w5204;
assign w5217 = ~w5215 & w5216;
assign w5218 = ~w5201 & ~w5202;
assign w5219 = ~w5217 & w5218;
assign w5220 = ~w5200 & ~w5219;
assign w5221 = ~w5199 & ~w5220;
assign w5222 = ~w5198 & ~w5221;
assign w5223 = ~w5197 & ~w5222;
assign w5224 = ~w5196 & ~w5223;
assign w5225 = ~pi135 & pi167;
assign w5226 = pi135 & ~pi167;
assign w5227 = pi136 & ~pi168;
assign w5228 = ~pi136 & pi168;
assign w5229 = ~pi137 & pi169;
assign w5230 = pi137 & ~pi169;
assign w5231 = pi138 & ~pi170;
assign w5232 = pi139 & ~pi171;
assign w5233 = pi140 & ~pi172;
assign w5234 = ~pi141 & pi173;
assign w5235 = pi141 & ~pi173;
assign w5236 = pi142 & ~pi174;
assign w5237 = ~w5235 & ~w5236;
assign w5238 = ~pi140 & pi172;
assign w5239 = ~w5234 & ~w5238;
assign w5240 = ~w5237 & w5239;
assign w5241 = ~w5232 & ~w5233;
assign w5242 = ~w5240 & w5241;
assign w5243 = ~pi138 & pi170;
assign w5244 = ~pi139 & pi171;
assign w5245 = ~w5243 & ~w5244;
assign w5246 = ~w5242 & w5245;
assign w5247 = ~w5230 & ~w5231;
assign w5248 = ~w5246 & w5247;
assign w5249 = ~w5228 & ~w5229;
assign w5250 = ~w5248 & w5249;
assign w5251 = ~w5226 & ~w5227;
assign w5252 = ~w5250 & w5251;
assign w5253 = ~w5225 & ~w5252;
assign w5254 = ~pi135 & pi191;
assign w5255 = pi135 & ~pi191;
assign w5256 = ~pi136 & pi192;
assign w5257 = pi136 & ~pi192;
assign w5258 = ~pi137 & pi193;
assign w5259 = pi137 & ~pi193;
assign w5260 = pi138 & ~pi194;
assign w5261 = ~pi139 & pi195;
assign w5262 = ~pi138 & pi194;
assign w5263 = pi139 & ~pi195;
assign w5264 = pi140 & ~pi196;
assign w5265 = ~pi140 & pi196;
assign w5266 = pi141 & ~pi197;
assign w5267 = ~pi141 & pi197;
assign w5268 = pi142 & ~pi198;
assign w5269 = ~w5267 & w5268;
assign w5270 = ~w5266 & ~w5269;
assign w5271 = ~w5265 & ~w5270;
assign w5272 = ~w5263 & ~w5264;
assign w5273 = ~w5271 & w5272;
assign w5274 = ~w5261 & ~w5262;
assign w5275 = ~w5273 & w5274;
assign w5276 = ~w5259 & ~w5260;
assign w5277 = ~w5275 & w5276;
assign w5278 = ~w5258 & ~w5277;
assign w5279 = ~w5257 & ~w5278;
assign w5280 = ~w5256 & ~w5279;
assign w5281 = ~w5255 & ~w5280;
assign w5282 = ~w5254 & ~w5281;
assign w5283 = ~w5253 & ~w5282;
assign w5284 = ~pi135 & pi151;
assign w5285 = pi136 & ~pi152;
assign w5286 = pi135 & ~pi151;
assign w5287 = pi137 & ~pi153;
assign w5288 = pi138 & ~pi154;
assign w5289 = ~pi138 & pi154;
assign w5290 = ~pi139 & pi155;
assign w5291 = pi139 & ~pi155;
assign w5292 = pi140 & ~pi156;
assign w5293 = ~pi141 & pi157;
assign w5294 = pi141 & ~pi157;
assign w5295 = pi142 & ~pi158;
assign w5296 = ~w5294 & ~w5295;
assign w5297 = ~pi140 & pi156;
assign w5298 = ~w5293 & ~w5297;
assign w5299 = ~w5296 & w5298;
assign w5300 = ~w5291 & ~w5292;
assign w5301 = ~w5299 & w5300;
assign w5302 = ~w5289 & ~w5290;
assign w5303 = ~w5301 & w5302;
assign w5304 = ~w5287 & ~w5288;
assign w5305 = ~w5303 & w5304;
assign w5306 = ~pi136 & pi152;
assign w5307 = ~pi137 & pi153;
assign w5308 = ~w5306 & ~w5307;
assign w5309 = ~w5305 & w5308;
assign w5310 = ~w5285 & ~w5286;
assign w5311 = ~w5309 & w5310;
assign w5312 = ~w5284 & ~w5311;
assign w5313 = ~pi135 & pi175;
assign w5314 = pi135 & ~pi175;
assign w5315 = ~pi136 & pi176;
assign w5316 = pi136 & ~pi176;
assign w5317 = ~pi137 & pi177;
assign w5318 = pi137 & ~pi177;
assign w5319 = pi138 & ~pi178;
assign w5320 = ~pi139 & pi179;
assign w5321 = ~pi138 & pi178;
assign w5322 = pi139 & ~pi179;
assign w5323 = pi140 & ~pi180;
assign w5324 = ~pi140 & pi180;
assign w5325 = pi141 & ~pi181;
assign w5326 = ~pi141 & pi181;
assign w5327 = pi142 & ~pi182;
assign w5328 = ~w5326 & w5327;
assign w5329 = ~w5325 & ~w5328;
assign w5330 = ~w5324 & ~w5329;
assign w5331 = ~w5322 & ~w5323;
assign w5332 = ~w5330 & w5331;
assign w5333 = ~w5320 & ~w5321;
assign w5334 = ~w5332 & w5333;
assign w5335 = ~w5318 & ~w5319;
assign w5336 = ~w5334 & w5335;
assign w5337 = ~w5317 & ~w5336;
assign w5338 = ~w5316 & ~w5337;
assign w5339 = ~w5315 & ~w5338;
assign w5340 = ~w5314 & ~w5339;
assign w5341 = ~w5313 & ~w5340;
assign w5342 = ~w5224 & ~w5312;
assign w5343 = ~w5341 & w5342;
assign w5344 = w5283 & w5343;
assign w5345 = w5195 & w5344;
assign w5346 = pi087 & w4714;
assign w5347 = pi135 & ~w5346;
assign w5348 = ~w1198 & w4707;
assign w5349 = ~pi135 & pi143;
assign w5350 = pi135 & ~pi143;
assign w5351 = pi136 & ~pi144;
assign w5352 = ~pi137 & pi145;
assign w5353 = ~pi136 & pi144;
assign w5354 = pi137 & ~pi145;
assign w5355 = pi138 & ~pi146;
assign w5356 = ~pi138 & pi146;
assign w5357 = ~pi139 & pi147;
assign w5358 = pi141 & ~pi149;
assign w5359 = ~pi141 & pi149;
assign w5360 = pi142 & ~pi150;
assign w5361 = ~w5359 & w5360;
assign w5362 = ~w5358 & ~w5361;
assign w5363 = ~pi148 & ~w5362;
assign w5364 = pi139 & ~pi147;
assign w5365 = pi148 & w5362;
assign w5366 = pi140 & ~w5365;
assign w5367 = ~w5363 & ~w5364;
assign w5368 = ~w5366 & w5367;
assign w5369 = ~w5356 & ~w5357;
assign w5370 = ~w5368 & w5369;
assign w5371 = ~w5354 & ~w5355;
assign w5372 = ~w5370 & w5371;
assign w5373 = ~w5352 & ~w5353;
assign w5374 = ~w5372 & w5373;
assign w5375 = ~w5350 & ~w5351;
assign w5376 = ~w5374 & w5375;
assign w5377 = ~w5349 & ~w5376;
assign w5378 = w4055 & ~w4715;
assign w5379 = ~w4725 & w5378;
assign w5380 = w2594 & ~w5347;
assign w5381 = w5379 & w5380;
assign w5382 = ~w950 & w5381;
assign w5383 = ~w1042 & ~w2532;
assign w5384 = ~w4711 & w5383;
assign w5385 = w5382 & w5384;
assign w5386 = ~w1948 & ~w3195;
assign w5387 = ~w3713 & w5386;
assign w5388 = w4060 & w5385;
assign w5389 = w5387 & w5388;
assign w5390 = w4063 & ~w4133;
assign w5391 = ~w4312 & w4721;
assign w5392 = w5390 & w5391;
assign w5393 = ~w5377 & w5389;
assign w5394 = w5392 & w5393;
assign w5395 = w5348 & w5394;
assign w5396 = w5345 & w5395;
assign w5397 = ~w28 & w4731;
assign w5398 = w2549 & w5397;
assign w5399 = ~w1014 & ~w2231;
assign w5400 = w2595 & w5399;
assign w5401 = w4723 & w5400;
assign w5402 = w5398 & w5401;
assign w5403 = ~w913 & w5402;
assign w5404 = ~w4054 & w5403;
assign w5405 = w852 & w5404;
assign w5406 = w5396 & w5405;
assign w5407 = ~w1921 & w5406;
assign w5408 = pi013 & w5407;
assign w5409 = (w4691 & w16251) | (w4691 & ~w4765) | (w16251 & ~w4765);
assign w5410 = (w4773 & ~w4827) | (w4773 & w16252) | (~w4827 & w16252);
assign w5411 = (w4769 & ~w4792) | (w4769 & w17552) | (~w4792 & w17552);
assign w5412 = (w4770 & ~w4792) | (w4770 & w17553) | (~w4792 & w17553);
assign w5413 = (~w4071 & ~w4781) | (~w4071 & w17030) | (~w4781 & w17030);
assign w5414 = (w4771 & ~w4755) | (w4771 & w17554) | (~w4755 & w17554);
assign w5415 = (w4777 & ~w4852) | (w4777 & w17555) | (~w4852 & w17555);
assign w5416 = ~w4705 & w4775;
assign w5417 = ~w5409 & ~w5410;
assign w5418 = w5413 & ~w5414;
assign w5419 = ~w5415 & ~w5416;
assign w5420 = w5418 & w5419;
assign w5421 = ~w5412 & w5417;
assign w5422 = w5420 & w5421;
assign w5423 = pi010 & w5422;
assign w5424 = ~w3949 & ~w4051;
assign w5425 = ~w4705 & w4750;
assign w5426 = (w4751 & ~w4827) | (w4751 & w16253) | (~w4827 & w16253);
assign w5427 = w4744 & ~w4854;
assign w5428 = ~w5425 & ~w5426;
assign w5429 = ~w5427 & w5428;
assign w5430 = (w4009 & ~w4686) | (w4009 & w17031) | (~w4686 & w17031);
assign w5431 = (~w3352 & ~w4096) | (~w3352 & w17556) | (~w4096 & w17556);
assign w5432 = (w4096 & w17557) | (w4096 & w17558) | (w17557 & w17558);
assign w5433 = (w4752 & ~w4792) | (w4752 & w17032) | (~w4792 & w17032);
assign w5434 = (w4745 & ~w4781) | (w4745 & w17033) | (~w4781 & w17033);
assign w5435 = w3978 & ~w4742;
assign w5436 = w3745 & ~w5435;
assign w5437 = (w5436 & ~w4755) | (w5436 & w17559) | (~w4755 & w17559);
assign w5438 = ~w5409 & w5437;
assign w5439 = ~w5430 & w5432;
assign w5440 = ~w5433 & ~w5434;
assign w5441 = w5439 & w5440;
assign w5442 = w5438 & w5441;
assign w5443 = ~w5425 & w17560;
assign w5444 = w5442 & w5443;
assign w5445 = pi009 & w5444;
assign w5446 = (w4104 & ~w4827) | (w4104 & w17034) | (~w4827 & w17034);
assign w5447 = (w4105 & ~w4755) | (w4105 & w17035) | (~w4755 & w17035);
assign w5448 = w4674 & ~w4705;
assign w5449 = (w4676 & ~w4852) | (w4676 & w17036) | (~w4852 & w17036);
assign w5450 = (w4679 & ~w4792) | (w4679 & w17037) | (~w4792 & w17037);
assign w5451 = w4313 & ~w4741;
assign w5452 = w4284 & ~w5451;
assign w5453 = (w5452 & ~w4686) | (w5452 & w17038) | (~w4686 & w17038);
assign w5454 = ~w5431 & w5453;
assign w5455 = ~w5413 & ~w5446;
assign w5456 = ~w5447 & ~w5448;
assign w5457 = ~w5449 & ~w5450;
assign w5458 = w5456 & w5457;
assign w5459 = w5454 & w5455;
assign w5460 = w5458 & w5459;
assign w5461 = w4672 & w5460;
assign w5462 = pi011 & w5461;
assign w5463 = (~w4051 & ~w4755) | (~w4051 & w18022) | (~w4755 & w18022);
assign w5464 = ~w4757 & w16256;
assign w5465 = ~w2291 & w4769;
assign w5466 = (w5465 & ~w4792) | (w5465 & w17039) | (~w4792 & w17039);
assign w5467 = w3048 & w4774;
assign w5468 = ~w4705 & w5467;
assign w5469 = ~w5466 & ~w5468;
assign w5470 = ~w5464 & w5469;
assign w5471 = ~w4094 & w17561;
assign w5472 = (w5471 & ~w4827) | (w5471 & w17040) | (~w4827 & w17040);
assign w5473 = (~w4163 & ~w4686) | (~w4163 & w17041) | (~w4686 & w17041);
assign w5474 = ~w5472 & ~w5473;
assign w5475 = (w3350 & ~w3419) | (w3350 & w17562) | (~w3419 & w17562);
assign w5476 = ~w883 & w5475;
assign w5477 = (w5476 & ~w4852) | (w5476 & w17563) | (~w4852 & w17563);
assign w5478 = w4742 & w5377;
assign w5479 = (w4852 & w17564) | (w4852 & w17565) | (w17564 & w17565);
assign w5480 = w5474 & w5479;
assign w5481 = w5470 & w5480;
assign w5482 = pi014 & w5481;
assign w5483 = ~w852 & w5475;
assign w5484 = (w5483 & ~w4852) | (w5483 & w17042) | (~w4852 & w17042);
assign w5485 = (~w4313 & ~w4686) | (~w4313 & w17043) | (~w4686 & w17043);
assign w5486 = ~w3387 & w17566;
assign w5487 = (w5486 & ~w4792) | (w5486 & w17044) | (~w4792 & w17044);
assign w5488 = w4071 & ~w4742;
assign w5489 = (~w5488 & ~w4781) | (~w5488 & w17045) | (~w4781 & w17045);
assign w5490 = w1261 & w4103;
assign w5491 = (w5490 & ~w4827) | (w5490 & w17046) | (~w4827 & w17046);
assign w5492 = ~w3978 & ~w4051;
assign w5493 = (w5492 & ~w4755) | (w5492 & w17047) | (~w4755 & w17047);
assign w5494 = ~w2990 & w4774;
assign w5495 = ~w4705 & w5494;
assign w5496 = ~w5409 & ~w5484;
assign w5497 = ~w5485 & ~w5487;
assign w5498 = ~w5489 & ~w5491;
assign w5499 = ~w5493 & ~w5495;
assign w5500 = w5498 & w5499;
assign w5501 = w5496 & w5497;
assign w5502 = w5500 & w5501;
assign w5503 = pi012 & w5502;
assign w5504 = (w4692 & ~w4765) | (w4692 & w16258) | (~w4765 & w16258);
assign w5505 = (~w2753 & ~w4686) | (~w2753 & w17048) | (~w4686 & w17048);
assign w5506 = (w4696 & ~w4852) | (w4696 & w17049) | (~w4852 & w17049);
assign w5507 = (w4689 & ~w4827) | (w4689 & w16259) | (~w4827 & w16259);
assign w5508 = (w4695 & ~w4755) | (w4695 & w17050) | (~w4755 & w17050);
assign w5509 = w2990 & ~w4742;
assign w5510 = (w4690 & ~w4792) | (w4690 & w17051) | (~w4792 & w17051);
assign w5511 = (w4698 & ~w4781) | (w4698 & w17052) | (~w4781 & w17052);
assign w5512 = w2724 & w3049;
assign w5513 = ~w5509 & w5512;
assign w5514 = (w4096 & w17567) | (w4096 & w17568) | (w17567 & w17568);
assign w5515 = ~w5504 & w5514;
assign w5516 = ~w5505 & ~w5506;
assign w5517 = ~w5507 & ~w5508;
assign w5518 = ~w5510 & ~w5511;
assign w5519 = w5517 & w5518;
assign w5520 = w5515 & w5516;
assign w5521 = w5519 & w5520;
assign w5522 = ~w4705 & w4774;
assign w5523 = ~w4705 & w17053;
assign w5524 = w2844 & w3169;
assign w5525 = ~w3254 & w5524;
assign w5526 = w2932 & ~w3225;
assign w5527 = ~w2961 & w5526;
assign w5528 = w5525 & w5527;
assign w5529 = ~w2873 & w5528;
assign w5530 = ~w4705 & w17569;
assign w5531 = w5521 & w5530;
assign w5532 = pi007 & w5531;
assign w5533 = w5409 & ~w5431;
assign w5534 = (w4759 & ~w4852) | (w4759 & w17054) | (~w4852 & w17054);
assign w5535 = (w4762 & ~w4827) | (w4762 & w16261) | (~w4827 & w16261);
assign w5536 = (w4761 & ~w4792) | (w4761 & w17055) | (~w4792 & w17055);
assign w5537 = ~w4705 & w4760;
assign w5538 = ~w5534 & ~w5535;
assign w5539 = ~w5536 & ~w5537;
assign w5540 = w5538 & w5539;
assign w5541 = w5533 & w5540;
assign w5542 = w2167 & ~w4797;
assign w5543 = w1920 & ~w2198;
assign w5544 = w5542 & w5543;
assign w5545 = (w4786 & ~w4827) | (w4786 & w16262) | (~w4827 & w16262);
assign w5546 = (w2473 & ~w4686) | (w2473 & w17056) | (~w4686 & w17056);
assign w5547 = ~w5545 & ~w5546;
assign w5548 = ~w4705 & w4787;
assign w5549 = (w4793 & ~w4755) | (w4793 & w17057) | (~w4755 & w17057);
assign w5550 = (w4788 & ~w4765) | (w4788 & w16263) | (~w4765 & w16263);
assign w5551 = (w4794 & ~w4781) | (w4794 & w17058) | (~w4781 & w17058);
assign w5552 = (w4789 & ~w4852) | (w4789 & w17059) | (~w4852 & w17059);
assign w5553 = ~w5549 & ~w5550;
assign w5554 = ~w5551 & ~w5552;
assign w5555 = w5553 & w5554;
assign w5556 = ~w2229 & ~w4742;
assign w5557 = w4796 & ~w5556;
assign w5558 = ~w3346 & w5557;
assign w5559 = w5411 & w5558;
assign w5560 = ~w5548 & w5559;
assign w5561 = w5547 & w5560;
assign w5562 = w5555 & w5561;
assign w5563 = w5544 & w5562;
assign w5564 = w4785 & w5563;
assign w5565 = pi003 & w1756;
assign w5566 = w4813 & ~w4831;
assign w5567 = ~w4705 & w4823;
assign w5568 = w3356 & ~w3420;
assign w5569 = (w5568 & ~w4852) | (w5568 & w17060) | (~w4852 & w17060);
assign w5570 = ~w5567 & ~w5569;
assign w5571 = (w1292 & ~w4685) | (w1292 & w17061) | (~w4685 & w17061);
assign w5572 = ~w1261 & ~w4742;
assign w5573 = (w4812 & ~w4755) | (w4812 & w17062) | (~w4755 & w17062);
assign w5574 = (w4811 & ~w4765) | (w4811 & w16264) | (~w4765 & w16264);
assign w5575 = (w4814 & ~w4781) | (w4814 & w17063) | (~w4781 & w17063);
assign w5576 = w4816 & ~w5572;
assign w5577 = w4102 & w17064;
assign w5578 = ~w4827 & w5577;
assign w5579 = ~w5571 & w5578;
assign w5580 = ~w5573 & w5579;
assign w5581 = ~w5574 & ~w5575;
assign w5582 = w5580 & w5581;
assign w5583 = ~w5566 & w5570;
assign w5584 = w5582 & w5583;
assign w5585 = w5565 & w5584;
assign w5586 = ~w1949 & w5558;
assign w5587 = w4769 & w5586;
assign w5588 = w5544 & w5587;
assign w5589 = ~w4831 & w5588;
assign w5590 = ~w5548 & w5589;
assign w5591 = w5547 & w5590;
assign w5592 = w5555 & w5591;
assign w5593 = w852 & ~w4742;
assign w5594 = ~w3337 & ~w3346;
assign w5595 = ~w4854 & w5594;
assign w5596 = (w16265 & ~w4852) | (w16265 & w17065) | (~w4852 & w17065);
assign w5597 = ~w5593 & w5596;
assign w5598 = (~w754 & ~w4686) | (~w754 & w17066) | (~w4686 & w17066);
assign w5599 = ~w4705 & w4845;
assign w5600 = (w4834 & ~w4781) | (w4834 & w17067) | (~w4781 & w17067);
assign w5601 = (w4846 & ~w4827) | (w4846 & w16266) | (~w4827 & w16266);
assign w5602 = (w4833 & ~w4755) | (w4833 & w17068) | (~w4755 & w17068);
assign w5603 = (w4832 & ~w4792) | (w4832 & w17570) | (~w4792 & w17570);
assign w5604 = ~w4765 & w4844;
assign w5605 = ~w5598 & ~w5604;
assign w5606 = ~w5599 & ~w5600;
assign w5607 = ~w5601 & ~w5602;
assign w5608 = ~w5603 & w5607;
assign w5609 = w5605 & w5606;
assign w5610 = w5608 & w5609;
assign w5611 = w5596 & w17571;
assign w5612 = w5609 & w17069;
assign w5613 = pi001 & w5612;
assign w5614 = ~w5585 & ~w5592;
assign w5615 = ~w5613 & w5614;
assign w5616 = ~w5564 & ~w5615;
assign w5617 = ~w5532 & ~w5541;
assign w5618 = ~w5616 & w5617;
assign w5619 = ~pi008 & w5541;
assign w5620 = ~w5444 & ~w5619;
assign w5621 = ~w5618 & w5620;
assign w5622 = ~w5408 & ~w5423;
assign w5623 = ~w5482 & ~w5503;
assign w5624 = w5622 & w5623;
assign w5625 = ~w5445 & ~w5462;
assign w5626 = w5624 & w5625;
assign w5627 = ~w5621 & w5626;
assign w5628 = (w5468 & ~w5521) | (w5468 & w16267) | (~w5521 & w16267);
assign w5629 = ~w5377 & ~w5407;
assign w5630 = (~w5629 & ~w5470) | (~w5629 & w17070) | (~w5470 & w17070);
assign w5631 = (w5466 & ~w5591) | (w5466 & w17071) | (~w5591 & w17071);
assign w5632 = (~w5458 & w17572) | (~w5458 & w17573) | (w17572 & w17573);
assign w5633 = ~w4163 & w5632;
assign w5634 = w5630 & ~w5631;
assign w5635 = ~w5628 & w5634;
assign w5636 = ~w5633 & w5635;
assign w5637 = (w5464 & ~w5442) | (w5464 & w16269) | (~w5442 & w16269);
assign w5638 = (~w4742 & ~w5500) | (~w4742 & w17072) | (~w5500 & w17072);
assign w5639 = (w1756 & w4831) | (w1756 & w16270) | (w4831 & w16270);
assign w5640 = w5570 & w5639;
assign w5641 = w5582 & w5640;
assign w5642 = w5472 & ~w5641;
assign w5643 = ~w5642 & w17574;
assign w5644 = ~w4854 & w5475;
assign w5645 = (w5644 & w16271) | (w5644 & ~w5610) | (w16271 & ~w5610);
assign w5646 = ~w883 & w5645;
assign w5647 = w5643 & ~w5646;
assign w5648 = w5636 & w5647;
assign w5649 = pi014 & w5648;
assign w5650 = w5474 & ~w5477;
assign w5651 = w5470 & w5650;
assign w5652 = ~pi151 & pi207;
assign w5653 = pi152 & ~pi208;
assign w5654 = pi151 & ~pi207;
assign w5655 = ~pi152 & pi208;
assign w5656 = ~pi153 & pi209;
assign w5657 = pi153 & ~pi209;
assign w5658 = pi154 & ~pi210;
assign w5659 = ~pi155 & pi211;
assign w5660 = ~pi154 & pi210;
assign w5661 = pi157 & ~pi213;
assign w5662 = ~pi157 & pi213;
assign w5663 = pi158 & ~pi214;
assign w5664 = ~w5662 & w5663;
assign w5665 = ~w5661 & ~w5664;
assign w5666 = ~pi212 & ~w5665;
assign w5667 = pi155 & ~pi211;
assign w5668 = pi212 & w5665;
assign w5669 = pi156 & ~w5668;
assign w5670 = ~w5666 & ~w5667;
assign w5671 = ~w5669 & w5670;
assign w5672 = ~w5659 & ~w5660;
assign w5673 = ~w5671 & w5672;
assign w5674 = ~w5657 & ~w5658;
assign w5675 = ~w5673 & w5674;
assign w5676 = ~w5655 & ~w5656;
assign w5677 = ~w5675 & w5676;
assign w5678 = ~w5653 & ~w5654;
assign w5679 = ~w5677 & w5678;
assign w5680 = ~w5652 & ~w5679;
assign w5681 = ~pi151 & pi223;
assign w5682 = pi151 & ~pi223;
assign w5683 = pi152 & ~pi224;
assign w5684 = ~pi153 & pi225;
assign w5685 = ~pi152 & pi224;
assign w5686 = pi153 & ~pi225;
assign w5687 = pi154 & ~pi226;
assign w5688 = ~pi154 & pi226;
assign w5689 = ~pi155 & pi227;
assign w5690 = pi157 & ~pi229;
assign w5691 = ~pi157 & pi229;
assign w5692 = pi158 & ~pi230;
assign w5693 = ~w5691 & w5692;
assign w5694 = ~w5690 & ~w5693;
assign w5695 = ~pi228 & ~w5694;
assign w5696 = pi155 & ~pi227;
assign w5697 = pi228 & w5694;
assign w5698 = pi156 & ~w5697;
assign w5699 = ~w5695 & ~w5696;
assign w5700 = ~w5698 & w5699;
assign w5701 = ~w5688 & ~w5689;
assign w5702 = ~w5700 & w5701;
assign w5703 = ~w5686 & ~w5687;
assign w5704 = ~w5702 & w5703;
assign w5705 = ~w5684 & ~w5685;
assign w5706 = ~w5704 & w5705;
assign w5707 = ~w5682 & ~w5683;
assign w5708 = ~w5706 & w5707;
assign w5709 = ~w5681 & ~w5708;
assign w5710 = ~pi151 & pi199;
assign w5711 = pi151 & ~pi199;
assign w5712 = pi152 & ~pi200;
assign w5713 = pi153 & ~pi201;
assign w5714 = pi154 & ~pi202;
assign w5715 = ~pi154 & pi202;
assign w5716 = ~pi155 & pi203;
assign w5717 = pi155 & ~pi203;
assign w5718 = pi156 & ~pi204;
assign w5719 = ~pi157 & pi205;
assign w5720 = pi157 & ~pi205;
assign w5721 = pi158 & ~pi206;
assign w5722 = ~w5720 & ~w5721;
assign w5723 = ~pi156 & pi204;
assign w5724 = ~w5719 & ~w5723;
assign w5725 = ~w5722 & w5724;
assign w5726 = ~w5717 & ~w5718;
assign w5727 = ~w5725 & w5726;
assign w5728 = ~w5715 & ~w5716;
assign w5729 = ~w5727 & w5728;
assign w5730 = ~w5713 & ~w5714;
assign w5731 = ~w5729 & w5730;
assign w5732 = ~pi152 & pi200;
assign w5733 = ~pi153 & pi201;
assign w5734 = ~w5732 & ~w5733;
assign w5735 = ~w5731 & w5734;
assign w5736 = ~w5711 & ~w5712;
assign w5737 = ~w5735 & w5736;
assign w5738 = ~w5710 & ~w5737;
assign w5739 = ~w5709 & ~w5738;
assign w5740 = ~w5680 & w5739;
assign w5741 = pi151 & ~pi191;
assign w5742 = ~pi151 & pi191;
assign w5743 = pi152 & ~pi192;
assign w5744 = ~pi152 & pi192;
assign w5745 = pi153 & ~pi193;
assign w5746 = ~pi153 & pi193;
assign w5747 = pi154 & ~pi194;
assign w5748 = ~pi154 & pi194;
assign w5749 = pi155 & ~pi195;
assign w5750 = ~pi155 & pi195;
assign w5751 = ~pi156 & pi196;
assign w5752 = pi157 & ~pi197;
assign w5753 = ~pi157 & pi197;
assign w5754 = pi158 & ~pi198;
assign w5755 = ~w5753 & w5754;
assign w5756 = ~w5752 & ~w5755;
assign w5757 = ~w5751 & ~w5756;
assign w5758 = pi156 & ~pi196;
assign w5759 = ~w5757 & ~w5758;
assign w5760 = ~w5750 & ~w5759;
assign w5761 = ~w5749 & ~w5760;
assign w5762 = ~w5748 & ~w5761;
assign w5763 = ~w5747 & ~w5762;
assign w5764 = ~w5746 & ~w5763;
assign w5765 = ~w5745 & ~w5764;
assign w5766 = ~w5744 & ~w5765;
assign w5767 = ~w5743 & ~w5766;
assign w5768 = ~w5742 & ~w5767;
assign w5769 = ~w5741 & ~w5768;
assign w5770 = w5740 & w5769;
assign w5771 = ~pi151 & pi167;
assign w5772 = pi152 & ~pi168;
assign w5773 = pi151 & ~pi167;
assign w5774 = ~pi153 & pi169;
assign w5775 = ~pi152 & pi168;
assign w5776 = ~pi154 & pi170;
assign w5777 = ~pi155 & pi171;
assign w5778 = pi157 & ~pi173;
assign w5779 = ~pi157 & pi173;
assign w5780 = pi158 & ~pi174;
assign w5781 = ~w5779 & w5780;
assign w5782 = ~w5778 & ~w5781;
assign w5783 = ~pi172 & ~w5782;
assign w5784 = pi155 & ~pi171;
assign w5785 = pi172 & w5782;
assign w5786 = pi156 & ~w5785;
assign w5787 = ~w5783 & ~w5784;
assign w5788 = ~w5786 & w5787;
assign w5789 = ~w5776 & ~w5777;
assign w5790 = ~w5788 & w5789;
assign w5791 = pi153 & ~pi169;
assign w5792 = pi154 & ~pi170;
assign w5793 = ~w5791 & ~w5792;
assign w5794 = ~w5790 & w5793;
assign w5795 = ~w5774 & ~w5775;
assign w5796 = ~w5794 & w5795;
assign w5797 = ~w5772 & ~w5773;
assign w5798 = ~w5796 & w5797;
assign w5799 = ~w5771 & ~w5798;
assign w5800 = ~pi151 & pi183;
assign w5801 = pi151 & ~pi183;
assign w5802 = pi152 & ~pi184;
assign w5803 = ~pi152 & pi184;
assign w5804 = ~pi153 & pi185;
assign w5805 = pi153 & ~pi185;
assign w5806 = pi154 & ~pi186;
assign w5807 = pi155 & ~pi187;
assign w5808 = pi156 & ~pi188;
assign w5809 = ~pi157 & pi189;
assign w5810 = pi157 & ~pi189;
assign w5811 = pi158 & ~pi190;
assign w5812 = ~w5810 & ~w5811;
assign w5813 = ~pi156 & pi188;
assign w5814 = ~w5809 & ~w5813;
assign w5815 = ~w5812 & w5814;
assign w5816 = ~w5807 & ~w5808;
assign w5817 = ~w5815 & w5816;
assign w5818 = ~pi154 & pi186;
assign w5819 = ~pi155 & pi187;
assign w5820 = ~w5818 & ~w5819;
assign w5821 = ~w5817 & w5820;
assign w5822 = ~w5805 & ~w5806;
assign w5823 = ~w5821 & w5822;
assign w5824 = ~w5803 & ~w5804;
assign w5825 = ~w5823 & w5824;
assign w5826 = ~w5801 & ~w5802;
assign w5827 = ~w5825 & w5826;
assign w5828 = ~w5800 & ~w5827;
assign w5829 = ~pi151 & pi175;
assign w5830 = pi151 & ~pi175;
assign w5831 = ~pi152 & pi176;
assign w5832 = pi152 & ~pi176;
assign w5833 = ~pi153 & pi177;
assign w5834 = pi153 & ~pi177;
assign w5835 = pi154 & ~pi178;
assign w5836 = ~pi154 & pi178;
assign w5837 = ~pi155 & pi179;
assign w5838 = pi157 & ~pi181;
assign w5839 = ~pi157 & pi181;
assign w5840 = pi158 & ~pi182;
assign w5841 = ~w5839 & w5840;
assign w5842 = ~w5838 & ~w5841;
assign w5843 = ~pi180 & ~w5842;
assign w5844 = pi155 & ~pi179;
assign w5845 = pi180 & w5842;
assign w5846 = pi156 & ~w5845;
assign w5847 = ~w5843 & ~w5844;
assign w5848 = ~w5846 & w5847;
assign w5849 = ~w5836 & ~w5837;
assign w5850 = ~w5848 & w5849;
assign w5851 = ~w5834 & ~w5835;
assign w5852 = ~w5850 & w5851;
assign w5853 = ~w5833 & ~w5852;
assign w5854 = ~w5832 & ~w5853;
assign w5855 = ~w5831 & ~w5854;
assign w5856 = ~w5830 & ~w5855;
assign w5857 = ~w5829 & ~w5856;
assign w5858 = ~w5799 & ~w5828;
assign w5859 = ~w5857 & w5858;
assign w5860 = w5770 & w5859;
assign w5861 = ~pi151 & pi271;
assign w5862 = pi151 & ~pi271;
assign w5863 = pi152 & ~pi272;
assign w5864 = pi153 & ~pi273;
assign w5865 = pi154 & ~pi274;
assign w5866 = ~pi154 & pi274;
assign w5867 = ~pi155 & pi275;
assign w5868 = pi155 & ~pi275;
assign w5869 = pi156 & ~pi276;
assign w5870 = ~pi157 & pi277;
assign w5871 = pi157 & ~pi277;
assign w5872 = pi158 & ~pi278;
assign w5873 = ~w5871 & ~w5872;
assign w5874 = ~pi156 & pi276;
assign w5875 = ~w5870 & ~w5874;
assign w5876 = ~w5873 & w5875;
assign w5877 = ~w5868 & ~w5869;
assign w5878 = ~w5876 & w5877;
assign w5879 = ~w5866 & ~w5867;
assign w5880 = ~w5878 & w5879;
assign w5881 = ~w5864 & ~w5865;
assign w5882 = ~w5880 & w5881;
assign w5883 = ~pi152 & pi272;
assign w5884 = ~pi153 & pi273;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = ~w5882 & w5885;
assign w5887 = ~w5862 & ~w5863;
assign w5888 = ~w5886 & w5887;
assign w5889 = ~w5861 & ~w5888;
assign w5890 = ~pi151 & pi255;
assign w5891 = pi152 & ~pi256;
assign w5892 = pi151 & ~pi255;
assign w5893 = ~pi152 & pi256;
assign w5894 = ~pi153 & pi257;
assign w5895 = pi153 & ~pi257;
assign w5896 = pi154 & ~pi258;
assign w5897 = ~pi154 & pi258;
assign w5898 = ~pi155 & pi259;
assign w5899 = pi155 & ~pi259;
assign w5900 = pi156 & ~pi260;
assign w5901 = ~pi157 & pi261;
assign w5902 = pi157 & ~pi261;
assign w5903 = pi158 & ~pi262;
assign w5904 = ~w5902 & ~w5903;
assign w5905 = ~pi156 & pi260;
assign w5906 = ~w5901 & ~w5905;
assign w5907 = ~w5904 & w5906;
assign w5908 = ~w5899 & ~w5900;
assign w5909 = ~w5907 & w5908;
assign w5910 = ~w5897 & ~w5898;
assign w5911 = ~w5909 & w5910;
assign w5912 = ~w5895 & ~w5896;
assign w5913 = ~w5911 & w5912;
assign w5914 = ~w5893 & ~w5894;
assign w5915 = ~w5913 & w5914;
assign w5916 = ~w5891 & ~w5892;
assign w5917 = ~w5915 & w5916;
assign w5918 = ~w5890 & ~w5917;
assign w5919 = ~pi151 & pi231;
assign w5920 = pi151 & ~pi231;
assign w5921 = pi152 & ~pi232;
assign w5922 = ~pi153 & pi233;
assign w5923 = ~pi152 & pi232;
assign w5924 = pi153 & ~pi233;
assign w5925 = pi154 & ~pi234;
assign w5926 = ~pi154 & pi234;
assign w5927 = ~pi155 & pi235;
assign w5928 = pi157 & ~pi237;
assign w5929 = ~pi157 & pi237;
assign w5930 = pi158 & ~pi238;
assign w5931 = ~w5929 & w5930;
assign w5932 = ~w5928 & ~w5931;
assign w5933 = ~pi236 & ~w5932;
assign w5934 = pi155 & ~pi235;
assign w5935 = pi236 & w5932;
assign w5936 = pi156 & ~w5935;
assign w5937 = ~w5933 & ~w5934;
assign w5938 = ~w5936 & w5937;
assign w5939 = ~w5926 & ~w5927;
assign w5940 = ~w5938 & w5939;
assign w5941 = ~w5924 & ~w5925;
assign w5942 = ~w5940 & w5941;
assign w5943 = ~w5922 & ~w5923;
assign w5944 = ~w5942 & w5943;
assign w5945 = ~w5920 & ~w5921;
assign w5946 = ~w5944 & w5945;
assign w5947 = ~w5919 & ~w5946;
assign w5948 = ~w5918 & ~w5947;
assign w5949 = ~w5889 & w5948;
assign w5950 = ~pi151 & pi239;
assign w5951 = pi151 & ~pi239;
assign w5952 = pi152 & ~pi240;
assign w5953 = ~pi153 & pi241;
assign w5954 = ~pi152 & pi240;
assign w5955 = pi153 & ~pi241;
assign w5956 = pi154 & ~pi242;
assign w5957 = ~pi154 & pi242;
assign w5958 = ~pi155 & pi243;
assign w5959 = pi157 & ~pi245;
assign w5960 = ~pi157 & pi245;
assign w5961 = pi158 & ~pi246;
assign w5962 = ~w5960 & w5961;
assign w5963 = ~w5959 & ~w5962;
assign w5964 = ~pi244 & ~w5963;
assign w5965 = pi155 & ~pi243;
assign w5966 = pi244 & w5963;
assign w5967 = pi156 & ~w5966;
assign w5968 = ~w5964 & ~w5965;
assign w5969 = ~w5967 & w5968;
assign w5970 = ~w5957 & ~w5958;
assign w5971 = ~w5969 & w5970;
assign w5972 = ~w5955 & ~w5956;
assign w5973 = ~w5971 & w5972;
assign w5974 = ~w5953 & ~w5954;
assign w5975 = ~w5973 & w5974;
assign w5976 = ~w5951 & ~w5952;
assign w5977 = ~w5975 & w5976;
assign w5978 = ~w5950 & ~w5977;
assign w5979 = ~pi151 & pi263;
assign w5980 = pi152 & ~pi264;
assign w5981 = pi151 & ~pi263;
assign w5982 = ~pi152 & pi264;
assign w5983 = ~pi153 & pi265;
assign w5984 = pi153 & ~pi265;
assign w5985 = pi154 & ~pi266;
assign w5986 = ~pi155 & pi267;
assign w5987 = ~pi154 & pi266;
assign w5988 = pi157 & ~pi269;
assign w5989 = ~pi157 & pi269;
assign w5990 = pi158 & ~pi270;
assign w5991 = ~w5989 & w5990;
assign w5992 = ~w5988 & ~w5991;
assign w5993 = ~pi268 & ~w5992;
assign w5994 = pi155 & ~pi267;
assign w5995 = pi268 & w5992;
assign w5996 = pi156 & ~w5995;
assign w5997 = ~w5993 & ~w5994;
assign w5998 = ~w5996 & w5997;
assign w5999 = ~w5986 & ~w5987;
assign w6000 = ~w5998 & w5999;
assign w6001 = ~w5984 & ~w5985;
assign w6002 = ~w6000 & w6001;
assign w6003 = ~w5982 & ~w5983;
assign w6004 = ~w6002 & w6003;
assign w6005 = ~w5980 & ~w5981;
assign w6006 = ~w6004 & w6005;
assign w6007 = ~w5979 & ~w6006;
assign w6008 = ~pi151 & pi247;
assign w6009 = pi151 & ~pi247;
assign w6010 = pi152 & ~pi248;
assign w6011 = ~pi152 & pi248;
assign w6012 = ~pi153 & pi249;
assign w6013 = pi153 & ~pi249;
assign w6014 = pi154 & ~pi250;
assign w6015 = pi155 & ~pi251;
assign w6016 = pi156 & ~pi252;
assign w6017 = ~pi157 & pi253;
assign w6018 = pi157 & ~pi253;
assign w6019 = pi158 & ~pi254;
assign w6020 = ~w6018 & ~w6019;
assign w6021 = ~pi156 & pi252;
assign w6022 = ~w6017 & ~w6021;
assign w6023 = ~w6020 & w6022;
assign w6024 = ~w6015 & ~w6016;
assign w6025 = ~w6023 & w6024;
assign w6026 = ~pi154 & pi250;
assign w6027 = ~pi155 & pi251;
assign w6028 = ~w6026 & ~w6027;
assign w6029 = ~w6025 & w6028;
assign w6030 = ~w6013 & ~w6014;
assign w6031 = ~w6029 & w6030;
assign w6032 = ~w6011 & ~w6012;
assign w6033 = ~w6031 & w6032;
assign w6034 = ~w6009 & ~w6010;
assign w6035 = ~w6033 & w6034;
assign w6036 = ~w6008 & ~w6035;
assign w6037 = ~w6007 & ~w6036;
assign w6038 = ~pi151 & pi215;
assign w6039 = pi151 & ~pi215;
assign w6040 = pi152 & ~pi216;
assign w6041 = ~pi152 & pi216;
assign w6042 = ~pi153 & pi217;
assign w6043 = pi153 & ~pi217;
assign w6044 = pi154 & ~pi218;
assign w6045 = pi155 & ~pi219;
assign w6046 = pi156 & ~pi220;
assign w6047 = ~pi157 & pi221;
assign w6048 = pi157 & ~pi221;
assign w6049 = pi158 & ~pi222;
assign w6050 = ~w6048 & ~w6049;
assign w6051 = ~pi156 & pi220;
assign w6052 = ~w6047 & ~w6051;
assign w6053 = ~w6050 & w6052;
assign w6054 = ~w6045 & ~w6046;
assign w6055 = ~w6053 & w6054;
assign w6056 = ~pi154 & pi218;
assign w6057 = ~pi155 & pi219;
assign w6058 = ~w6056 & ~w6057;
assign w6059 = ~w6055 & w6058;
assign w6060 = ~w6043 & ~w6044;
assign w6061 = ~w6059 & w6060;
assign w6062 = ~w6041 & ~w6042;
assign w6063 = ~w6061 & w6062;
assign w6064 = ~w6039 & ~w6040;
assign w6065 = ~w6063 & w6064;
assign w6066 = ~w6038 & ~w6065;
assign w6067 = ~w5978 & ~w6066;
assign w6068 = w6037 & w6067;
assign w6069 = w5949 & w6068;
assign w6070 = ~pi151 & pi159;
assign w6071 = pi152 & ~pi160;
assign w6072 = pi151 & ~pi159;
assign w6073 = pi153 & ~pi161;
assign w6074 = pi154 & ~pi162;
assign w6075 = pi155 & ~pi163;
assign w6076 = pi156 & ~pi164;
assign w6077 = ~pi157 & pi165;
assign w6078 = pi157 & ~pi165;
assign w6079 = pi158 & ~pi166;
assign w6080 = ~w6078 & ~w6079;
assign w6081 = ~pi156 & pi164;
assign w6082 = ~w6077 & ~w6081;
assign w6083 = ~w6080 & w6082;
assign w6084 = ~w6075 & ~w6076;
assign w6085 = ~w6083 & w6084;
assign w6086 = ~pi154 & pi162;
assign w6087 = ~pi155 & pi163;
assign w6088 = ~w6086 & ~w6087;
assign w6089 = ~w6085 & w6088;
assign w6090 = ~w6073 & ~w6074;
assign w6091 = ~w6089 & w6090;
assign w6092 = ~pi152 & pi160;
assign w6093 = ~pi153 & pi161;
assign w6094 = ~w6092 & ~w6093;
assign w6095 = ~w6091 & w6094;
assign w6096 = ~w6071 & ~w6072;
assign w6097 = ~w6095 & w6096;
assign w6098 = ~w6070 & ~w6097;
assign w6099 = ~w27 & w4717;
assign w6100 = w4062 & w4720;
assign w6101 = w6099 & w6100;
assign w6102 = w2627 & w4712;
assign w6103 = ~w4312 & ~w5376;
assign w6104 = w4707 & w6103;
assign w6105 = w4708 & w6104;
assign w6106 = w6102 & w6105;
assign w6107 = pi039 & pi055;
assign w6108 = pi071 & w6107;
assign w6109 = pi135 & w6108;
assign w6110 = w5346 & w6109;
assign w6111 = pi151 & ~w6110;
assign w6112 = ~w4715 & ~w5349;
assign w6113 = w5397 & w6112;
assign w6114 = w4735 & w6113;
assign w6115 = w1327 & ~w6111;
assign w6116 = ~w2162 & w6115;
assign w6117 = ~w787 & w6116;
assign w6118 = ~w2872 & ~w5311;
assign w6119 = w6117 & w6118;
assign w6120 = ~w6098 & w6119;
assign w6121 = ~w3653 & w6114;
assign w6122 = w6120 & w6121;
assign w6123 = w6101 & w6122;
assign w6124 = w6069 & w6123;
assign w6125 = w6106 & w6124;
assign w6126 = w5860 & w6125;
assign w6127 = w5651 & w6126;
assign w6128 = w5470 & w17073;
assign w6129 = pi015 & w6128;
assign w6130 = w4519 & w5632;
assign w6131 = ~w4705 & w17575;
assign w6132 = (w6131 & ~w5521) | (w6131 & w16273) | (~w5521 & w16273);
assign w6133 = ~w2444 & w5411;
assign w6134 = (w6133 & ~w5591) | (w6133 & w17074) | (~w5591 & w17074);
assign w6135 = ~w5224 & ~w5407;
assign w6136 = w5470 & w17075;
assign w6137 = ~w6134 & w6136;
assign w6138 = ~w6132 & w6137;
assign w6139 = ~w6130 & w6138;
assign w6140 = ~w3683 & w5463;
assign w6141 = (w6140 & ~w5442) | (w6140 & w16274) | (~w5442 & w16274);
assign w6142 = w691 & w5644;
assign w6143 = (w6142 & ~w5610) | (w6142 & w16275) | (~w5610 & w16275);
assign w6144 = w4103 & ~w4828;
assign w6145 = ~w5641 & w6144;
assign w6146 = ~w5641 & w16276;
assign w6147 = ~w6143 & ~w6146;
assign w6148 = ~w6141 & w6147;
assign w6149 = w6139 & w6148;
assign w6150 = w5478 & w6098;
assign w6151 = w6149 & w6150;
assign w6152 = pi016 & w6151;
assign w6153 = ~w3714 & w5463;
assign w6154 = (w6153 & ~w5442) | (w6153 & w16277) | (~w5442 & w16277);
assign w6155 = (w5523 & ~w5521) | (w5523 & w16278) | (~w5521 & w16278);
assign w6156 = ~w5641 & w16279;
assign w6157 = ~w4134 & ~w4687;
assign w6158 = (w6157 & w16280) | (w6157 & ~w5460) | (w16280 & ~w5460);
assign w6159 = w5411 & ~w5592;
assign w6160 = (w16281 & ~w5591) | (w16281 & w17076) | (~w5591 & w17076);
assign w6161 = w913 & w5644;
assign w6162 = (w6161 & ~w5610) | (w6161 & w16282) | (~w5610 & w16282);
assign w6163 = (w5470 & w17077) | (w5470 & w17078) | (w17077 & w17078);
assign w6164 = ~w5638 & w6163;
assign w6165 = ~w6154 & ~w6155;
assign w6166 = ~w6156 & ~w6158;
assign w6167 = ~w6160 & ~w6162;
assign w6168 = w6166 & w6167;
assign w6169 = w6164 & w6165;
assign w6170 = w6168 & w6169;
assign w6171 = ~pi013 & w6170;
assign w6172 = (w5599 & ~w5521) | (w5599 & w16283) | (~w5521 & w16283);
assign w6173 = (w883 & ~w5470) | (w883 & w17079) | (~w5470 & w17079);
assign w6174 = (w5463 & ~w5442) | (w5463 & w16284) | (~w5442 & w16284);
assign w6175 = w278 & w6174;
assign w6176 = ~w5612 & ~w6173;
assign w6177 = ~w6172 & w6176;
assign w6178 = ~w6175 & w6177;
assign w6179 = (w5598 & ~w5460) | (w5598 & w16285) | (~w5460 & w16285);
assign w6180 = (w5604 & ~w5540) | (w5604 & w16286) | (~w5540 & w16286);
assign w6181 = ~w913 & ~w5407;
assign w6182 = w4837 & ~w6181;
assign w6183 = w5596 & w6182;
assign w6184 = (w5593 & ~w5500) | (w5593 & w17080) | (~w5500 & w17080);
assign w6185 = w5601 & ~w5641;
assign w6186 = (w5600 & ~w5420) | (w5600 & w16287) | (~w5420 & w16287);
assign w6187 = (w5603 & ~w5591) | (w5603 & w17081) | (~w5591 & w17081);
assign w6188 = ~w6184 & ~w6185;
assign w6189 = ~w6186 & ~w6187;
assign w6190 = w6188 & w6189;
assign w6191 = w822 & w6183;
assign w6192 = ~w6180 & w6191;
assign w6193 = ~w6179 & w6192;
assign w6194 = w6190 & w6193;
assign w6195 = w6178 & w6194;
assign w6196 = pi001 & w6195;
assign w6197 = (w5508 & ~w5442) | (w5508 & w16288) | (~w5442 & w16288);
assign w6198 = (~w5609 & w17082) | (~w5609 & w17083) | (w17082 & w17083);
assign w6199 = (~w5458 & w17084) | (~w5458 & w17085) | (w17084 & w17085);
assign w6200 = w3019 & ~w5431;
assign w6201 = ~w2723 & w6200;
assign w6202 = (w6201 & w5540) | (w6201 & w16291) | (w5540 & w16291);
assign w6203 = (w5509 & ~w5500) | (w5509 & w17086) | (~w5500 & w17086);
assign w6204 = (w5511 & ~w5420) | (w5511 & w16292) | (~w5420 & w16292);
assign w6205 = (~w3048 & ~w5470) | (~w3048 & w17087) | (~w5470 & w17087);
assign w6206 = (w5510 & ~w5591) | (w5510 & w17088) | (~w5591 & w17088);
assign w6207 = w5507 & ~w5641;
assign w6208 = w3197 & ~w5407;
assign w6209 = (w5540 & w17576) | (w5540 & w17577) | (w17576 & w17577);
assign w6210 = ~w6203 & ~w6204;
assign w6211 = ~w6205 & ~w6206;
assign w6212 = ~w6207 & w6211;
assign w6213 = w6209 & w6210;
assign w6214 = w6132 & ~w6197;
assign w6215 = ~w6198 & ~w6199;
assign w6216 = w6214 & w6215;
assign w6217 = w6212 & w6213;
assign w6218 = w6216 & w6217;
assign w6219 = w6217 & w16293;
assign w6220 = pi007 & w6219;
assign w6221 = (~w5609 & w17578) | (~w5609 & w17579) | (w17578 & w17579);
assign w6222 = (w5413 & ~w5420) | (w5413 & w16295) | (~w5420 & w16295);
assign w6223 = (w5412 & ~w5591) | (w5412 & w17089) | (~w5591 & w17089);
assign w6224 = (w5414 & ~w5442) | (w5414 & w16296) | (~w5442 & w16296);
assign w6225 = (w5409 & ~w5540) | (w5409 & w16297) | (~w5540 & w16297);
assign w6226 = w5410 & ~w5641;
assign w6227 = w6222 & ~w6223;
assign w6228 = ~w6225 & ~w6226;
assign w6229 = w6227 & w6228;
assign w6230 = ~w6221 & ~w6224;
assign w6231 = w6228 & w17580;
assign w6232 = (w5522 & ~w5521) | (w5522 & w17581) | (~w5521 & w17581);
assign w6233 = ~w3287 & w6232;
assign w6234 = w6231 & ~w6233;
assign w6235 = pi010 & w6234;
assign w6236 = (w5549 & ~w5442) | (w5549 & w16298) | (~w5442 & w16298);
assign w6237 = (~w5609 & w17090) | (~w5609 & w17091) | (w17090 & w17091);
assign w6238 = ~w6236 & ~w6237;
assign w6239 = (~w5458 & w17092) | (~w5458 & w17093) | (w17092 & w17093);
assign w6240 = (~w4831 & ~w5591) | (~w4831 & w17582) | (~w5591 & w17582);
assign w6241 = (w5548 & ~w5521) | (w5548 & w16301) | (~w5521 & w16301);
assign w6242 = w5545 & ~w5641;
assign w6243 = (w2291 & ~w5470) | (w2291 & w17094) | (~w5470 & w17094);
assign w6244 = (~w5539 & w18118) | (~w5539 & w18119) | (w18118 & w18119);
assign w6245 = (w5551 & ~w5420) | (w5551 & w16303) | (~w5420 & w16303);
assign w6246 = ~w6244 & ~w6245;
assign w6247 = (w5556 & ~w5500) | (w5556 & w17095) | (~w5500 & w17095);
assign w6248 = ~w2540 & ~w3387;
assign w6249 = w1949 & ~w5406;
assign w6250 = w4795 & ~w6249;
assign w6251 = w5542 & w6250;
assign w6252 = w6248 & w6251;
assign w6253 = (w6252 & w5641) | (w6252 & w16304) | (w5641 & w16304);
assign w6254 = ~w6243 & ~w6247;
assign w6255 = w6253 & w6254;
assign w6256 = ~w6241 & w6246;
assign w6257 = w6255 & w6256;
assign w6258 = w3376 & w5543;
assign w6259 = (w16305 & ~w5591) | (w16305 & w17096) | (~w5591 & w17096);
assign w6260 = ~w6239 & w6259;
assign w6261 = w6238 & w6260;
assign w6262 = w6257 & w6261;
assign w6263 = pi005 & w6262;
assign w6264 = (~w5610 & w17097) | (~w5610 & w17098) | (w17097 & w17098);
assign w6265 = (w5536 & ~w5591) | (w5536 & w17099) | (~w5591 & w17099);
assign w6266 = (w5537 & ~w5521) | (w5537 & w18023) | (~w5521 & w18023);
assign w6267 = w5535 & ~w5641;
assign w6268 = (w5533 & ~w5539) | (w5533 & w18024) | (~w5539 & w18024);
assign w6269 = ~w6265 & w6268;
assign w6270 = ~w6267 & w6269;
assign w6271 = ~w6266 & w6270;
assign w6272 = w6270 & w16306;
assign w6273 = pi008 & w6272;
assign w6274 = (w5448 & ~w5521) | (w5448 & w16307) | (~w5521 & w16307);
assign w6275 = w4134 & ~w5407;
assign w6276 = w4282 & ~w4687;
assign w6277 = (w5451 & ~w5500) | (w5451 & w17100) | (~w5500 & w17100);
assign w6278 = w5446 & ~w5641;
assign w6279 = (w4163 & ~w5470) | (w4163 & w17101) | (~w5470 & w17101);
assign w6280 = (w5450 & ~w5591) | (w5450 & w17102) | (~w5591 & w17102);
assign w6281 = ~w6275 & w6276;
assign w6282 = (w5420 & w18025) | (w5420 & w18026) | (w18025 & w18026);
assign w6283 = ~w6277 & ~w6278;
assign w6284 = ~w6279 & ~w6280;
assign w6285 = w6283 & w6284;
assign w6286 = ~w6274 & w6282;
assign w6287 = w6283 & w18027;
assign w6288 = (w5447 & ~w5442) | (w5447 & w16308) | (~w5442 & w16308);
assign w6289 = (~w5458 & w17103) | (~w5458 & w17104) | (w17103 & w17104);
assign w6290 = ~w6288 & w6289;
assign w6291 = (~w5609 & w17105) | (~w5609 & w17106) | (w17105 & w17106);
assign w6292 = w4672 & ~w6291;
assign w6293 = w6290 & w6292;
assign w6294 = w6285 & w17583;
assign w6295 = pi011 & w6294;
assign w6296 = (~w5458 & w17107) | (~w5458 & w17108) | (w17107 & w17108);
assign w6297 = w5491 & ~w5641;
assign w6298 = ~w6222 & ~w6297;
assign w6299 = ~w6297 & w17584;
assign w6300 = (w5487 & ~w5591) | (w5487 & w17109) | (~w5591 & w17109);
assign w6301 = (w5495 & ~w5521) | (w5495 & w16312) | (~w5521 & w16312);
assign w6302 = (w5493 & ~w5442) | (w5493 & w16313) | (~w5442 & w16313);
assign w6303 = w5484 & ~w5612;
assign w6304 = ~w6301 & ~w6302;
assign w6305 = ~w6303 & w6304;
assign w6306 = w6298 & w16314;
assign w6307 = w6305 & w6306;
assign w6308 = w6306 & w17110;
assign w6309 = pi012 & w6308;
assign w6310 = w3362 & ~w4828;
assign w6311 = (w1104 & ~w5470) | (w1104 & w18321) | (~w5470 & w18321);
assign w6312 = w1043 & ~w5407;
assign w6313 = ~w1388 & w6222;
assign w6314 = (w5572 & ~w5500) | (w5572 & w17111) | (~w5500 & w17111);
assign w6315 = (w5566 & ~w5591) | (w5566 & w17112) | (~w5591 & w17112);
assign w6316 = (w5567 & ~w5521) | (w5567 & w16315) | (~w5521 & w16315);
assign w6317 = (w5574 & ~w5540) | (w5574 & w16316) | (~w5540 & w16316);
assign w6318 = (w5540 & w17113) | (w5540 & w17114) | (w17113 & w17114);
assign w6319 = (~w5609 & w17115) | (~w5609 & w17116) | (w17115 & w17116);
assign w6320 = (~w5458 & w17117) | (~w5458 & w17118) | (w17117 & w17118);
assign w6321 = (w5573 & ~w5442) | (w5573 & w16319) | (~w5442 & w16319);
assign w6322 = w1359 & ~w6312;
assign w6323 = (w5470 & w17585) | (w5470 & w17586) | (w17585 & w17586);
assign w6324 = ~w6314 & ~w6315;
assign w6325 = w6323 & w6324;
assign w6326 = ~w6313 & ~w6316;
assign w6327 = w6318 & ~w6319;
assign w6328 = ~w6320 & ~w6321;
assign w6329 = w6327 & w6328;
assign w6330 = w6325 & w6326;
assign w6331 = w6329 & w6330;
assign w6332 = w6310 & w6331;
assign w6333 = w4102 & ~w5641;
assign w6334 = ~w1073 & w3310;
assign w6335 = w6333 & w6334;
assign w6336 = w3355 & w6335;
assign w6337 = w6332 & w6336;
assign w6338 = (w3743 & ~w5470) | (w3743 & w17119) | (~w5470 & w17119);
assign w6339 = w5426 & ~w5641;
assign w6340 = w3714 & ~w5407;
assign w6341 = (w5433 & ~w5591) | (w5433 & w17120) | (~w5591 & w17120);
assign w6342 = (w5435 & ~w5500) | (w5435 & w17121) | (~w5500 & w17121);
assign w6343 = ~w5422 & w5434;
assign w6344 = (~w5458 & w17122) | (~w5458 & w17123) | (w17122 & w17123);
assign w6345 = (w5425 & ~w5521) | (w5425 & w16322) | (~w5521 & w16322);
assign w6346 = (w5427 & ~w5610) | (w5427 & w16323) | (~w5610 & w16323);
assign w6347 = w3685 & ~w6340;
assign w6348 = w5432 & w6347;
assign w6349 = ~w6225 & w6348;
assign w6350 = ~w6338 & ~w6339;
assign w6351 = ~w6341 & ~w6342;
assign w6352 = ~w6343 & w6351;
assign w6353 = w6349 & w6350;
assign w6354 = w6174 & ~w6344;
assign w6355 = ~w6345 & ~w6346;
assign w6356 = w6354 & w6355;
assign w6357 = w6352 & w6353;
assign w6358 = w6356 & w6357;
assign w6359 = w6357 & w16324;
assign w6360 = pi009 & w6359;
assign w6361 = ~w6170 & ~w6196;
assign w6362 = ~w6235 & ~w6263;
assign w6363 = ~w6273 & ~w6295;
assign w6364 = w6362 & w6363;
assign w6365 = ~w6220 & w6361;
assign w6366 = ~w6309 & ~w6337;
assign w6367 = ~w6360 & w6366;
assign w6368 = w6364 & w6365;
assign w6369 = w6367 & w6368;
assign w6370 = ~w5648 & ~w6171;
assign w6371 = ~w6369 & w6370;
assign w6372 = ~w5649 & ~w6129;
assign w6373 = ~w6152 & w6372;
assign w6374 = ~w6371 & w6373;
assign w6375 = w6069 & ~w6128;
assign w6376 = pi015 & w6375;
assign w6377 = w1756 & ~w3346;
assign w6378 = ~w1073 & w4815;
assign w6379 = w6377 & w6378;
assign w6380 = ~w5641 & w17587;
assign w6381 = w6330 & w16325;
assign w6382 = w6145 & ~w6381;
assign w6383 = ~w1329 & w6382;
assign w6384 = w4062 & w6104;
assign w6385 = w4721 & w6098;
assign w6386 = w6099 & w6114;
assign w6387 = w6385 & w6386;
assign w6388 = w4713 & w6387;
assign w6389 = w6384 & w6388;
assign w6390 = (~w16274 & w17124) | (~w16274 & w17125) | (w17124 & w17125);
assign w6391 = w6147 & w6390;
assign w6392 = w6139 & w6391;
assign w6393 = (w6098 & ~w6139) | (w6098 & w16326) | (~w6139 & w16326);
assign w6394 = ~w4490 & w5632;
assign w6395 = (w6394 & ~w6287) | (w6394 & w16327) | (~w6287 & w16327);
assign w6396 = ~w5312 & ~w5407;
assign w6397 = (w6396 & ~w6168) | (w6396 & w17588) | (~w6168 & w17588);
assign w6398 = ~w789 & w5645;
assign w6399 = (w6398 & ~w6194) | (w6398 & w17126) | (~w6194 & w17126);
assign w6400 = ~w6393 & ~w6395;
assign w6401 = ~w6397 & ~w6399;
assign w6402 = w6400 & w6401;
assign w6403 = ~w6383 & w6402;
assign w6404 = ~w3654 & w6174;
assign w6405 = (w6404 & ~w6357) | (w6404 & w17589) | (~w6357 & w17589);
assign w6406 = (w6159 & ~w6257) | (w6159 & w16328) | (~w6257 & w16328);
assign w6407 = ~w2164 & w6406;
assign w6408 = w6217 & w16329;
assign w6409 = ~w2873 & w6232;
assign w6410 = ~w6408 & w6409;
assign w6411 = ~w6407 & ~w6410;
assign w6412 = (~w5481 & ~w5647) | (~w5481 & w17127) | (~w5647 & w17127);
assign w6413 = w5860 & ~w6412;
assign w6414 = ~w6405 & w6413;
assign w6415 = w6411 & w6414;
assign w6416 = w6403 & w6415;
assign w6417 = w6376 & w6416;
assign w6418 = (w6162 & ~w6194) | (w6162 & w17128) | (~w6194 & w17128);
assign w6419 = w5312 & ~w6128;
assign w6420 = w5195 & ~w5431;
assign w6421 = w6156 & ~w6381;
assign w6422 = w6155 & ~w6219;
assign w6423 = ~w5648 & w16330;
assign w6424 = (w5224 & ~w6139) | (w5224 & w16331) | (~w6139 & w16331);
assign w6425 = ~w5341 & ~w5407;
assign w6426 = (w6425 & ~w6168) | (w6425 & w17590) | (~w6168 & w17590);
assign w6427 = (w6154 & ~w6357) | (w6154 & w17591) | (~w6357 & w17591);
assign w6428 = (w6158 & ~w6287) | (w6158 & w16332) | (~w6287 & w16332);
assign w6429 = (w6160 & ~w6257) | (w6160 & w16333) | (~w6257 & w16333);
assign w6430 = w5283 & w6420;
assign w6431 = ~w6419 & w6430;
assign w6432 = w6306 & w17592;
assign w6433 = ~w6418 & w6432;
assign w6434 = ~w6424 & w6426;
assign w6435 = ~w6428 & ~w6429;
assign w6436 = w6434 & w6435;
assign w6437 = ~w6421 & w6433;
assign w6438 = ~w6422 & ~w6423;
assign w6439 = ~w6427 & w6438;
assign w6440 = w6436 & w6437;
assign w6441 = w6439 & w6440;
assign w6442 = ~pi013 & w6441;
assign w6443 = w5860 & w6375;
assign w6444 = (w5647 & w17129) | (w5647 & w17130) | (w17129 & w17130);
assign w6445 = ~w6405 & w6444;
assign w6446 = w6411 & w6445;
assign w6447 = w6403 & w6446;
assign w6448 = (w5629 & ~w6168) | (w5629 & w17593) | (~w6168 & w17593);
assign w6449 = (w5631 & ~w6257) | (w5631 & w16335) | (~w6257 & w16335);
assign w6450 = (w5632 & ~w6287) | (w5632 & w16336) | (~w6287 & w16336);
assign w6451 = (~w6287 & w5633) | (~w6287 & w17131) | (w5633 & w17131);
assign w6452 = (w5637 & ~w6357) | (w5637 & w17594) | (~w6357 & w17594);
assign w6453 = (w5646 & ~w6194) | (w5646 & w17132) | (~w6194 & w17132);
assign w6454 = w5642 & ~w6381;
assign w6455 = w5628 & ~w6219;
assign w6456 = ~w5648 & w16337;
assign w6457 = ~w6448 & ~w6449;
assign w6458 = ~w6453 & w6457;
assign w6459 = ~w6451 & w6456;
assign w6460 = ~w6452 & w17133;
assign w6461 = w6458 & w6459;
assign w6462 = w6460 & w6461;
assign w6463 = ~w6447 & ~w6462;
assign w6464 = w6225 & ~w6272;
assign w6465 = (w6343 & ~w6231) | (w6343 & w16338) | (~w6231 & w16338);
assign w6466 = ~w6464 & ~w6465;
assign w6467 = (~w5461 & ~w6287) | (~w5461 & w16339) | (~w6287 & w16339);
assign w6468 = (~w6287 & w17134) | (~w6287 & w17135) | (w17134 & w17135);
assign w6469 = ~w6219 & w6345;
assign w6470 = w3920 & ~w4757;
assign w6471 = ~w5444 & w6470;
assign w6472 = (w6471 & ~w6357) | (w6471 & w17595) | (~w6357 & w17595);
assign w6473 = (w6340 & ~w6168) | (w6340 & w18028) | (~w6168 & w18028);
assign w6474 = (w6342 & ~w6306) | (w6342 & w18029) | (~w6306 & w18029);
assign w6475 = (w6346 & ~w6194) | (w6346 & w17136) | (~w6194 & w17136);
assign w6476 = w3654 & ~w6128;
assign w6477 = w3625 & ~w5431;
assign w6478 = ~w6476 & w6477;
assign w6479 = ~w6473 & w6478;
assign w6480 = ~w6474 & ~w6475;
assign w6481 = w6479 & w6480;
assign w6482 = w6466 & ~w6468;
assign w6483 = ~w6469 & w6472;
assign w6484 = w6482 & w6483;
assign w6485 = w6481 & w6484;
assign w6486 = w6339 & ~w6381;
assign w6487 = w3743 & w6412;
assign w6488 = (w3683 & ~w6139) | (w3683 & w16340) | (~w6139 & w16340);
assign w6489 = (w6341 & ~w6257) | (w6341 & w16341) | (~w6257 & w16341);
assign w6490 = ~w6488 & ~w6489;
assign w6491 = ~w6486 & w6490;
assign w6492 = ~w6487 & w6491;
assign w6493 = w6491 & w17137;
assign w6494 = w6485 & w6493;
assign w6495 = pi009 & w6494;
assign w6496 = w6277 & ~w6308;
assign w6497 = (w6288 & ~w6357) | (w6288 & w17596) | (~w6357 & w17596);
assign w6498 = w6278 & ~w6381;
assign w6499 = ~w6219 & w6274;
assign w6500 = (~w6229 & w17138) | (~w6229 & w17139) | (w17138 & w17139);
assign w6501 = (w6279 & ~w5647) | (w6279 & w17140) | (~w5647 & w17140);
assign w6502 = (w6280 & ~w6257) | (w6280 & w16343) | (~w6257 & w16343);
assign w6503 = (~w4519 & ~w6139) | (~w4519 & w16344) | (~w6139 & w16344);
assign w6504 = (w6275 & ~w6168) | (w6275 & w17597) | (~w6168 & w17597);
assign w6505 = (w6291 & ~w6194) | (w6291 & w17598) | (~w6194 & w17598);
assign w6506 = w4490 & ~w6127;
assign w6507 = w4402 & ~w6506;
assign w6508 = ~w6500 & w6507;
assign w6509 = ~w6501 & ~w6502;
assign w6510 = ~w6503 & ~w6504;
assign w6511 = ~w6505 & w6510;
assign w6512 = w6508 & w6509;
assign w6513 = ~w6496 & ~w6497;
assign w6514 = ~w6498 & ~w6499;
assign w6515 = w6513 & w6514;
assign w6516 = w6511 & w6512;
assign w6517 = w6515 & w6516;
assign w6518 = w4461 & ~w5431;
assign w6519 = w4282 & w6518;
assign w6520 = (~w6287 & w17141) | (~w6287 & w17142) | (w17141 & w17142);
assign w6521 = w4670 & w6520;
assign w6522 = ~w4551 & w6521;
assign w6523 = w6516 & w16345;
assign w6524 = ~w6219 & w6233;
assign w6525 = (w6221 & ~w6194) | (w6221 & w17143) | (~w6194 & w17143);
assign w6526 = ~w6381 & w18030;
assign w6527 = (w6224 & ~w6357) | (w6224 & w17599) | (~w6357 & w17599);
assign w6528 = (w6223 & ~w6257) | (w6223 & w16346) | (~w6257 & w16346);
assign w6529 = ~w6464 & w6500;
assign w6530 = ~w6525 & ~w6528;
assign w6531 = w6529 & w6530;
assign w6532 = ~w6524 & ~w6527;
assign w6533 = w6531 & w16347;
assign w6534 = pi010 & w6533;
assign w6535 = w6207 & ~w6381;
assign w6536 = (w2695 & ~w6139) | (w2695 & w16348) | (~w6139 & w16348);
assign w6537 = (w6199 & ~w6287) | (w6199 & w16349) | (~w6287 & w16349);
assign w6538 = (w6208 & ~w6168) | (w6208 & w17600) | (~w6168 & w17600);
assign w6539 = (w6205 & ~w5647) | (w6205 & w17144) | (~w5647 & w17144);
assign w6540 = ~w6536 & ~w6537;
assign w6541 = ~w6538 & ~w6539;
assign w6542 = w6540 & w6541;
assign w6543 = (w6206 & ~w6257) | (w6206 & w16350) | (~w6257 & w16350);
assign w6544 = (w6204 & ~w6229) | (w6204 & w16351) | (~w6229 & w16351);
assign w6545 = (w2873 & ~w5470) | (w2873 & w18031) | (~w5470 & w18031);
assign w6546 = (w6197 & ~w6357) | (w6197 & w17601) | (~w6357 & w17601);
assign w6547 = (w6198 & ~w6194) | (w6198 & w17145) | (~w6194 & w17145);
assign w6548 = (w6203 & ~w6306) | (w6203 & w18032) | (~w6306 & w18032);
assign w6549 = w6202 & ~w6545;
assign w6550 = (w6229 & w17602) | (w6229 & w17603) | (w17602 & w17603);
assign w6551 = ~w6543 & w6550;
assign w6552 = ~w6547 & ~w6548;
assign w6553 = w6552 & w16352;
assign w6554 = w5528 & w6232;
assign w6555 = ~w6219 & w6554;
assign w6556 = ~w6535 & w6555;
assign w6557 = w6542 & w6556;
assign w6558 = w6553 & w6557;
assign w6559 = ~pi007 & w6558;
assign w6560 = w789 & ~w6128;
assign w6561 = w660 & ~w6560;
assign w6562 = ~w4854 & ~w6195;
assign w6563 = w2634 & ~w3420;
assign w6564 = ~w5612 & w6563;
assign w6565 = w4835 & w6564;
assign w6566 = w6562 & w6565;
assign w6567 = (~w6229 & w17146) | (~w6229 & w17147) | (w17146 & w17147);
assign w6568 = w6172 & ~w6219;
assign w6569 = (w6175 & ~w6357) | (w6175 & w17604) | (~w6357 & w17604);
assign w6570 = ~w6381 & w17605;
assign w6571 = (w6184 & ~w6306) | (w6184 & w17148) | (~w6306 & w17148);
assign w6572 = (w6173 & ~w5636) | (w6173 & w17606) | (~w5636 & w17606);
assign w6573 = ~w6567 & ~w6571;
assign w6574 = ~w6572 & w6573;
assign w6575 = ~w6568 & ~w6569;
assign w6576 = w6575 & w17149;
assign w6577 = (~w6287 & w17607) | (~w6287 & w17608) | (w17607 & w17608);
assign w6578 = (w6187 & ~w6257) | (w6187 & w16354) | (~w6257 & w16354);
assign w6579 = ~w691 & ~w6392;
assign w6580 = (~w5407 & ~w6168) | (~w5407 & w17609) | (~w6168 & w17609);
assign w6581 = (w6181 & ~w6168) | (w6181 & w18033) | (~w6168 & w18033);
assign w6582 = ~w6180 & ~w6578;
assign w6583 = ~w6579 & w6582;
assign w6584 = ~w6577 & ~w6581;
assign w6585 = w6583 & w6584;
assign w6586 = w6576 & w6585;
assign w6587 = w249 & ~w4847;
assign w6588 = ~w821 & w6587;
assign w6589 = pi001 & w5594;
assign w6590 = w6588 & w6589;
assign w6591 = w6561 & w6590;
assign w6592 = w6566 & w6591;
assign w6593 = w6586 & w6592;
assign w6594 = (w6236 & ~w6357) | (w6236 & w17610) | (~w6357 & w17610);
assign w6595 = (w6243 & ~w5647) | (w6243 & w17150) | (~w5647 & w17150);
assign w6596 = (~w6246 & ~w6231) | (~w6246 & w16355) | (~w6231 & w16355);
assign w6597 = (w6249 & ~w6168) | (w6249 & w17611) | (~w6168 & w17611);
assign w6598 = (w6239 & ~w6287) | (w6239 & w16356) | (~w6287 & w16356);
assign w6599 = (w2444 & ~w6139) | (w2444 & w16357) | (~w6139 & w16357);
assign w6600 = w6299 & w6305;
assign w6601 = w6247 & ~w6600;
assign w6602 = ~w6595 & ~w6596;
assign w6603 = ~w6597 & ~w6598;
assign w6604 = ~w6599 & ~w6601;
assign w6605 = w6603 & w6604;
assign w6606 = ~w6594 & w6602;
assign w6607 = w6605 & w6606;
assign w6608 = w6242 & ~w6381;
assign w6609 = (w6237 & ~w6194) | (w6237 & w17151) | (~w6194 & w17151);
assign w6610 = ~w6608 & ~w6609;
assign w6611 = w2164 & ~w6128;
assign w6612 = ~w2134 & w2322;
assign w6613 = w2416 & w6612;
assign w6614 = ~w4797 & w6613;
assign w6615 = (w6614 & w6128) | (w6614 & w17612) | (w6128 & w17612);
assign w6616 = ~w6241 & w6615;
assign w6617 = w5529 & w6615;
assign w6618 = (~w6616 & ~w6218) | (~w6616 & w16358) | (~w6218 & w16358);
assign w6619 = w6240 & w6248;
assign w6620 = (w6619 & ~w6257) | (w6619 & w16359) | (~w6257 & w16359);
assign w6621 = w2104 & ~w2198;
assign w6622 = w2043 & w6621;
assign w6623 = w1920 & w6622;
assign w6624 = w3376 & w6623;
assign w6625 = w6620 & w6624;
assign w6626 = ~w6618 & w6625;
assign w6627 = w6610 & w6626;
assign w6628 = w6607 & w6627;
assign w6629 = ~w6558 & ~w6628;
assign w6630 = w6310 & ~w6381;
assign w6631 = w1329 & ~w6128;
assign w6632 = (w6319 & ~w6194) | (w6319 & w18322) | (~w6194 & w18322);
assign w6633 = w1358 & ~w6392;
assign w6634 = w6318 & ~w6631;
assign w6635 = (w6194 & w17152) | (w6194 & w17153) | (w17152 & w17153);
assign w6636 = ~w6633 & w6635;
assign w6637 = (w6321 & ~w6357) | (w6321 & w17613) | (~w6357 & w17613);
assign w6638 = (w6314 & ~w6306) | (w6314 & w17614) | (~w6306 & w17614);
assign w6639 = (w6312 & ~w6168) | (w6312 & w17615) | (~w6168 & w17615);
assign w6640 = (w6313 & ~w6231) | (w6313 & w16361) | (~w6231 & w16361);
assign w6641 = (w6315 & ~w6257) | (w6315 & w16362) | (~w6257 & w16362);
assign w6642 = (w6320 & ~w6287) | (w6320 & w16363) | (~w6287 & w16363);
assign w6643 = (w6311 & ~w5647) | (w6311 & w17154) | (~w5647 & w17154);
assign w6644 = ~w6638 & ~w6639;
assign w6645 = ~w6640 & ~w6641;
assign w6646 = ~w6642 & ~w6643;
assign w6647 = w6645 & w6646;
assign w6648 = ~w6637 & w6644;
assign w6649 = w6647 & w6648;
assign w6650 = ~w6219 & w6316;
assign w6651 = w6630 & ~w6650;
assign w6652 = w6636 & w6651;
assign w6653 = w6649 & w6652;
assign w6654 = w6336 & w6653;
assign w6655 = w6629 & ~w6654;
assign w6656 = ~w6593 & w6655;
assign w6657 = w6610 & ~w6618;
assign w6658 = w6607 & w6657;
assign w6659 = w6622 & w6658;
assign w6660 = w3376 & ~w5592;
assign w6661 = w6248 & ~w6262;
assign w6662 = ~w4831 & w6661;
assign w6663 = w1920 & w6662;
assign w6664 = ~pi005 & w6663;
assign w6665 = w6660 & w6664;
assign w6666 = w6659 & w6665;
assign w6667 = ~w6494 & ~w6559;
assign w6668 = ~w6666 & w6667;
assign w6669 = ~w6656 & w6668;
assign w6670 = ~w6523 & ~w6534;
assign w6671 = ~w6495 & w6670;
assign w6672 = ~w6669 & w6671;
assign w6673 = (w6303 & ~w6194) | (w6303 & w17155) | (~w6194 & w17155);
assign w6674 = (w6300 & ~w6257) | (w6300 & w17616) | (~w6257 & w17616);
assign w6675 = ~w6219 & w6301;
assign w6676 = ~w6294 & w6296;
assign w6677 = w6297 & ~w6381;
assign w6678 = (w6302 & ~w6357) | (w6302 & w17617) | (~w6357 & w17617);
assign w6679 = ~w6307 & ~w6500;
assign w6680 = ~w6673 & ~w6674;
assign w6681 = ~w6676 & w6680;
assign w6682 = ~w6675 & w6679;
assign w6683 = ~w6677 & ~w6678;
assign w6684 = w6682 & w6683;
assign w6685 = w6681 & w6684;
assign w6686 = ~pi011 & w6523;
assign w6687 = ~w6685 & ~w6686;
assign w6688 = ~w6672 & w6687;
assign w6689 = pi012 & w6685;
assign w6690 = ~w6441 & ~w6689;
assign w6691 = ~w6688 & w6690;
assign w6692 = ~w6442 & w6463;
assign w6693 = ~w6691 & w6692;
assign w6694 = pi014 & w6462;
assign w6695 = ~w6097 & w6384;
assign w6696 = ~pi167 & pi255;
assign w6697 = pi168 & ~pi256;
assign w6698 = pi167 & ~pi255;
assign w6699 = ~pi168 & pi256;
assign w6700 = ~pi169 & pi257;
assign w6701 = pi169 & ~pi257;
assign w6702 = pi170 & ~pi258;
assign w6703 = ~pi170 & pi258;
assign w6704 = ~pi171 & pi259;
assign w6705 = pi173 & ~pi261;
assign w6706 = ~pi173 & pi261;
assign w6707 = pi174 & ~pi262;
assign w6708 = ~w6706 & w6707;
assign w6709 = ~w6705 & ~w6708;
assign w6710 = ~pi260 & ~w6709;
assign w6711 = pi171 & ~pi259;
assign w6712 = pi260 & w6709;
assign w6713 = pi172 & ~w6712;
assign w6714 = ~w6710 & ~w6711;
assign w6715 = ~w6713 & w6714;
assign w6716 = ~w6703 & ~w6704;
assign w6717 = ~w6715 & w6716;
assign w6718 = ~w6701 & ~w6702;
assign w6719 = ~w6717 & w6718;
assign w6720 = ~w6699 & ~w6700;
assign w6721 = ~w6719 & w6720;
assign w6722 = ~w6697 & ~w6698;
assign w6723 = ~w6721 & w6722;
assign w6724 = ~w6696 & ~w6723;
assign w6725 = ~pi167 & pi247;
assign w6726 = pi168 & ~pi248;
assign w6727 = pi167 & ~pi247;
assign w6728 = ~pi169 & pi249;
assign w6729 = ~pi168 & pi248;
assign w6730 = pi169 & ~pi249;
assign w6731 = pi170 & ~pi250;
assign w6732 = ~pi170 & pi250;
assign w6733 = ~pi171 & pi251;
assign w6734 = pi173 & ~pi253;
assign w6735 = ~pi173 & pi253;
assign w6736 = pi174 & ~pi254;
assign w6737 = ~w6735 & w6736;
assign w6738 = ~w6734 & ~w6737;
assign w6739 = ~pi252 & ~w6738;
assign w6740 = pi171 & ~pi251;
assign w6741 = pi252 & w6738;
assign w6742 = pi172 & ~w6741;
assign w6743 = ~w6739 & ~w6740;
assign w6744 = ~w6742 & w6743;
assign w6745 = ~w6732 & ~w6733;
assign w6746 = ~w6744 & w6745;
assign w6747 = ~w6730 & ~w6731;
assign w6748 = ~w6746 & w6747;
assign w6749 = ~w6728 & ~w6729;
assign w6750 = ~w6748 & w6749;
assign w6751 = ~w6726 & ~w6727;
assign w6752 = ~w6750 & w6751;
assign w6753 = ~w6725 & ~w6752;
assign w6754 = ~w6724 & ~w6753;
assign w6755 = ~pi167 & pi271;
assign w6756 = pi168 & ~pi272;
assign w6757 = pi167 & ~pi271;
assign w6758 = pi169 & ~pi273;
assign w6759 = pi170 & ~pi274;
assign w6760 = ~pi170 & pi274;
assign w6761 = ~pi171 & pi275;
assign w6762 = pi171 & ~pi275;
assign w6763 = pi172 & ~pi276;
assign w6764 = ~pi173 & pi277;
assign w6765 = pi173 & ~pi277;
assign w6766 = pi174 & ~pi278;
assign w6767 = ~w6765 & ~w6766;
assign w6768 = ~pi172 & pi276;
assign w6769 = ~w6764 & ~w6768;
assign w6770 = ~w6767 & w6769;
assign w6771 = ~w6762 & ~w6763;
assign w6772 = ~w6770 & w6771;
assign w6773 = ~w6760 & ~w6761;
assign w6774 = ~w6772 & w6773;
assign w6775 = ~w6758 & ~w6759;
assign w6776 = ~w6774 & w6775;
assign w6777 = ~pi168 & pi272;
assign w6778 = ~pi169 & pi273;
assign w6779 = ~w6777 & ~w6778;
assign w6780 = ~w6776 & w6779;
assign w6781 = ~w6756 & ~w6757;
assign w6782 = ~w6780 & w6781;
assign w6783 = ~w6755 & ~w6782;
assign w6784 = ~pi167 & pi263;
assign w6785 = pi167 & ~pi263;
assign w6786 = pi168 & ~pi264;
assign w6787 = ~pi168 & pi264;
assign w6788 = ~pi169 & pi265;
assign w6789 = pi169 & ~pi265;
assign w6790 = pi170 & ~pi266;
assign w6791 = pi171 & ~pi267;
assign w6792 = pi172 & ~pi268;
assign w6793 = ~pi173 & pi269;
assign w6794 = pi173 & ~pi269;
assign w6795 = pi174 & ~pi270;
assign w6796 = ~w6794 & ~w6795;
assign w6797 = ~pi172 & pi268;
assign w6798 = ~w6793 & ~w6797;
assign w6799 = ~w6796 & w6798;
assign w6800 = ~w6791 & ~w6792;
assign w6801 = ~w6799 & w6800;
assign w6802 = ~pi170 & pi266;
assign w6803 = ~pi171 & pi267;
assign w6804 = ~w6802 & ~w6803;
assign w6805 = ~w6801 & w6804;
assign w6806 = ~w6789 & ~w6790;
assign w6807 = ~w6805 & w6806;
assign w6808 = ~w6787 & ~w6788;
assign w6809 = ~w6807 & w6808;
assign w6810 = ~w6785 & ~w6786;
assign w6811 = ~w6809 & w6810;
assign w6812 = ~w6784 & ~w6811;
assign w6813 = ~w6783 & ~w6812;
assign w6814 = ~pi167 & pi239;
assign w6815 = pi167 & ~pi239;
assign w6816 = pi168 & ~pi240;
assign w6817 = ~pi168 & pi240;
assign w6818 = ~pi169 & pi241;
assign w6819 = pi169 & ~pi241;
assign w6820 = pi170 & ~pi242;
assign w6821 = ~pi171 & pi243;
assign w6822 = ~pi170 & pi242;
assign w6823 = pi173 & ~pi245;
assign w6824 = ~pi173 & pi245;
assign w6825 = pi174 & ~pi246;
assign w6826 = ~w6824 & w6825;
assign w6827 = ~w6823 & ~w6826;
assign w6828 = ~pi244 & ~w6827;
assign w6829 = pi171 & ~pi243;
assign w6830 = pi244 & w6827;
assign w6831 = pi172 & ~w6830;
assign w6832 = ~w6828 & ~w6829;
assign w6833 = ~w6831 & w6832;
assign w6834 = ~w6821 & ~w6822;
assign w6835 = ~w6833 & w6834;
assign w6836 = ~w6819 & ~w6820;
assign w6837 = ~w6835 & w6836;
assign w6838 = ~w6817 & ~w6818;
assign w6839 = ~w6837 & w6838;
assign w6840 = ~w6815 & ~w6816;
assign w6841 = ~w6839 & w6840;
assign w6842 = ~w6814 & ~w6841;
assign w6843 = ~pi167 & pi231;
assign w6844 = pi167 & ~pi231;
assign w6845 = pi168 & ~pi232;
assign w6846 = ~pi168 & pi232;
assign w6847 = ~pi169 & pi233;
assign w6848 = pi169 & ~pi233;
assign w6849 = pi170 & ~pi234;
assign w6850 = pi171 & ~pi235;
assign w6851 = pi172 & ~pi236;
assign w6852 = ~pi173 & pi237;
assign w6853 = pi173 & ~pi237;
assign w6854 = pi174 & ~pi238;
assign w6855 = ~w6853 & ~w6854;
assign w6856 = ~pi172 & pi236;
assign w6857 = ~w6852 & ~w6856;
assign w6858 = ~w6855 & w6857;
assign w6859 = ~w6850 & ~w6851;
assign w6860 = ~w6858 & w6859;
assign w6861 = ~pi170 & pi234;
assign w6862 = ~pi171 & pi235;
assign w6863 = ~w6861 & ~w6862;
assign w6864 = ~w6860 & w6863;
assign w6865 = ~w6848 & ~w6849;
assign w6866 = ~w6864 & w6865;
assign w6867 = ~w6846 & ~w6847;
assign w6868 = ~w6866 & w6867;
assign w6869 = ~w6844 & ~w6845;
assign w6870 = ~w6868 & w6869;
assign w6871 = ~w6843 & ~w6870;
assign w6872 = ~w6842 & ~w6871;
assign w6873 = ~pi167 & pi223;
assign w6874 = pi167 & ~pi223;
assign w6875 = pi168 & ~pi224;
assign w6876 = ~pi169 & pi225;
assign w6877 = ~pi168 & pi224;
assign w6878 = pi169 & ~pi225;
assign w6879 = pi170 & ~pi226;
assign w6880 = ~pi171 & pi227;
assign w6881 = ~pi170 & pi226;
assign w6882 = pi173 & ~pi229;
assign w6883 = ~pi173 & pi229;
assign w6884 = pi174 & ~pi230;
assign w6885 = ~w6883 & w6884;
assign w6886 = ~w6882 & ~w6885;
assign w6887 = ~pi228 & ~w6886;
assign w6888 = pi171 & ~pi227;
assign w6889 = pi228 & w6886;
assign w6890 = pi172 & ~w6889;
assign w6891 = ~w6887 & ~w6888;
assign w6892 = ~w6890 & w6891;
assign w6893 = ~w6880 & ~w6881;
assign w6894 = ~w6892 & w6893;
assign w6895 = ~w6878 & ~w6879;
assign w6896 = ~w6894 & w6895;
assign w6897 = ~w6876 & ~w6877;
assign w6898 = ~w6896 & w6897;
assign w6899 = ~w6874 & ~w6875;
assign w6900 = ~w6898 & w6899;
assign w6901 = ~w6873 & ~w6900;
assign w6902 = ~pi167 & pi215;
assign w6903 = pi168 & ~pi216;
assign w6904 = pi167 & ~pi215;
assign w6905 = pi169 & ~pi217;
assign w6906 = pi170 & ~pi218;
assign w6907 = ~pi170 & pi218;
assign w6908 = ~pi171 & pi219;
assign w6909 = pi171 & ~pi219;
assign w6910 = pi172 & ~pi220;
assign w6911 = ~pi173 & pi221;
assign w6912 = pi173 & ~pi221;
assign w6913 = pi174 & ~pi222;
assign w6914 = ~w6912 & ~w6913;
assign w6915 = ~pi172 & pi220;
assign w6916 = ~w6911 & ~w6915;
assign w6917 = ~w6914 & w6916;
assign w6918 = ~w6909 & ~w6910;
assign w6919 = ~w6917 & w6918;
assign w6920 = ~w6907 & ~w6908;
assign w6921 = ~w6919 & w6920;
assign w6922 = ~w6905 & ~w6906;
assign w6923 = ~w6921 & w6922;
assign w6924 = ~pi168 & pi216;
assign w6925 = ~pi169 & pi217;
assign w6926 = ~w6924 & ~w6925;
assign w6927 = ~w6923 & w6926;
assign w6928 = ~w6903 & ~w6904;
assign w6929 = ~w6927 & w6928;
assign w6930 = ~w6902 & ~w6929;
assign w6931 = w6813 & ~w6930;
assign w6932 = ~w6901 & w6931;
assign w6933 = w6754 & w6932;
assign w6934 = w6872 & w6933;
assign w6935 = ~pi167 & pi175;
assign w6936 = pi168 & ~pi176;
assign w6937 = pi167 & ~pi175;
assign w6938 = ~pi168 & pi176;
assign w6939 = ~pi169 & pi177;
assign w6940 = pi169 & ~pi177;
assign w6941 = pi170 & ~pi178;
assign w6942 = ~pi170 & pi178;
assign w6943 = ~pi171 & pi179;
assign w6944 = pi171 & ~pi179;
assign w6945 = pi172 & ~pi180;
assign w6946 = ~pi173 & pi181;
assign w6947 = pi173 & ~pi181;
assign w6948 = pi174 & ~pi182;
assign w6949 = ~w6947 & ~w6948;
assign w6950 = ~pi172 & pi180;
assign w6951 = ~w6946 & ~w6950;
assign w6952 = ~w6949 & w6951;
assign w6953 = ~w6944 & ~w6945;
assign w6954 = ~w6952 & w6953;
assign w6955 = ~w6942 & ~w6943;
assign w6956 = ~w6954 & w6955;
assign w6957 = ~w6940 & ~w6941;
assign w6958 = ~w6956 & w6957;
assign w6959 = ~w6938 & ~w6939;
assign w6960 = ~w6958 & w6959;
assign w6961 = ~w6936 & ~w6937;
assign w6962 = ~w6960 & w6961;
assign w6963 = ~w6935 & ~w6962;
assign w6964 = w2546 & w4712;
assign w6965 = w4720 & w6964;
assign w6966 = ~w616 & w620;
assign w6967 = ~w612 & w6966;
assign w6968 = w626 & ~w6967;
assign w6969 = w4056 & ~w6070;
assign w6970 = w6112 & w6969;
assign w6971 = ~pi167 & pi191;
assign w6972 = pi167 & ~pi191;
assign w6973 = ~pi168 & pi192;
assign w6974 = pi168 & ~pi192;
assign w6975 = ~pi169 & pi193;
assign w6976 = pi169 & ~pi193;
assign w6977 = pi170 & ~pi194;
assign w6978 = ~pi171 & pi195;
assign w6979 = ~pi170 & pi194;
assign w6980 = pi171 & ~pi195;
assign w6981 = pi172 & ~pi196;
assign w6982 = ~pi172 & pi196;
assign w6983 = pi173 & ~pi197;
assign w6984 = ~pi173 & pi197;
assign w6985 = pi174 & ~pi198;
assign w6986 = ~w6984 & w6985;
assign w6987 = ~w6983 & ~w6986;
assign w6988 = ~w6982 & ~w6987;
assign w6989 = ~w6980 & ~w6981;
assign w6990 = ~w6988 & w6989;
assign w6991 = ~w6978 & ~w6979;
assign w6992 = ~w6990 & w6991;
assign w6993 = ~w6976 & ~w6977;
assign w6994 = ~w6992 & w6993;
assign w6995 = ~w6975 & ~w6994;
assign w6996 = ~w6974 & ~w6995;
assign w6997 = ~w6973 & ~w6996;
assign w6998 = ~w6972 & ~w6997;
assign w6999 = ~w6971 & ~w6998;
assign w7000 = ~pi167 & pi207;
assign w7001 = pi168 & ~pi208;
assign w7002 = pi167 & ~pi207;
assign w7003 = ~pi169 & pi209;
assign w7004 = ~pi168 & pi208;
assign w7005 = ~pi170 & pi210;
assign w7006 = ~pi171 & pi211;
assign w7007 = pi173 & ~pi213;
assign w7008 = ~pi173 & pi213;
assign w7009 = pi174 & ~pi214;
assign w7010 = ~w7008 & w7009;
assign w7011 = ~w7007 & ~w7010;
assign w7012 = ~pi212 & ~w7011;
assign w7013 = pi171 & ~pi211;
assign w7014 = pi212 & w7011;
assign w7015 = pi172 & ~w7014;
assign w7016 = ~w7012 & ~w7013;
assign w7017 = ~w7015 & w7016;
assign w7018 = ~w7005 & ~w7006;
assign w7019 = ~w7017 & w7018;
assign w7020 = pi169 & ~pi209;
assign w7021 = pi170 & ~pi210;
assign w7022 = ~w7020 & ~w7021;
assign w7023 = ~w7019 & w7022;
assign w7024 = ~w7003 & ~w7004;
assign w7025 = ~w7023 & w7024;
assign w7026 = ~w7001 & ~w7002;
assign w7027 = ~w7025 & w7026;
assign w7028 = ~w7000 & ~w7027;
assign w7029 = ~pi167 & pi199;
assign w7030 = pi167 & ~pi199;
assign w7031 = pi168 & ~pi200;
assign w7032 = ~pi168 & pi200;
assign w7033 = ~pi169 & pi201;
assign w7034 = pi169 & ~pi201;
assign w7035 = pi170 & ~pi202;
assign w7036 = pi171 & ~pi203;
assign w7037 = pi172 & ~pi204;
assign w7038 = ~pi173 & pi205;
assign w7039 = pi173 & ~pi205;
assign w7040 = pi174 & ~pi206;
assign w7041 = ~w7039 & ~w7040;
assign w7042 = ~pi172 & pi204;
assign w7043 = ~w7038 & ~w7042;
assign w7044 = ~w7041 & w7043;
assign w7045 = ~w7036 & ~w7037;
assign w7046 = ~w7044 & w7045;
assign w7047 = ~pi170 & pi202;
assign w7048 = ~pi171 & pi203;
assign w7049 = ~w7047 & ~w7048;
assign w7050 = ~w7046 & w7049;
assign w7051 = ~w7034 & ~w7035;
assign w7052 = ~w7050 & w7051;
assign w7053 = ~w7032 & ~w7033;
assign w7054 = ~w7052 & w7053;
assign w7055 = ~w7030 & ~w7031;
assign w7056 = ~w7054 & w7055;
assign w7057 = ~w7029 & ~w7056;
assign w7058 = ~w7028 & ~w7057;
assign w7059 = ~pi167 & pi183;
assign w7060 = pi167 & ~pi183;
assign w7061 = pi168 & ~pi184;
assign w7062 = pi169 & ~pi185;
assign w7063 = pi170 & ~pi186;
assign w7064 = ~pi170 & pi186;
assign w7065 = ~pi171 & pi187;
assign w7066 = pi171 & ~pi187;
assign w7067 = pi172 & ~pi188;
assign w7068 = ~pi173 & pi189;
assign w7069 = pi173 & ~pi189;
assign w7070 = pi174 & ~pi190;
assign w7071 = ~w7069 & ~w7070;
assign w7072 = ~pi172 & pi188;
assign w7073 = ~w7068 & ~w7072;
assign w7074 = ~w7071 & w7073;
assign w7075 = ~w7066 & ~w7067;
assign w7076 = ~w7074 & w7075;
assign w7077 = ~w7064 & ~w7065;
assign w7078 = ~w7076 & w7077;
assign w7079 = ~w7062 & ~w7063;
assign w7080 = ~w7078 & w7079;
assign w7081 = ~pi168 & pi184;
assign w7082 = ~pi169 & pi185;
assign w7083 = ~w7081 & ~w7082;
assign w7084 = ~w7080 & w7083;
assign w7085 = ~w7060 & ~w7061;
assign w7086 = ~w7084 & w7085;
assign w7087 = ~w7059 & ~w7086;
assign w7088 = ~w6999 & ~w7087;
assign w7089 = w7058 & w7088;
assign w7090 = ~w1071 & w6970;
assign w7091 = ~w2132 & w4733;
assign w7092 = ~w6968 & w7091;
assign w7093 = w7090 & w7092;
assign w7094 = ~w2960 & ~w3594;
assign w7095 = ~w4341 & w4716;
assign w7096 = ~w5252 & w7095;
assign w7097 = w7093 & w7094;
assign w7098 = ~w6963 & w7097;
assign w7099 = ~w5798 & w7096;
assign w7100 = w6965 & w7099;
assign w7101 = w4061 & w7098;
assign w7102 = w7100 & w7101;
assign w7103 = w6695 & w7102;
assign w7104 = w6934 & w7089;
assign w7105 = w7103 & w7104;
assign w7106 = w6149 & w7105;
assign w7107 = pi151 & pi167;
assign w7108 = w5346 & w7107;
assign w7109 = w6109 & w7108;
assign w7110 = pi167 & ~w7109;
assign w7111 = ~w28 & w4728;
assign w7112 = ~w7110 & w7111;
assign w7113 = w6149 & w17618;
assign w7114 = pi017 & w7113;
assign w7115 = w6132 & ~w6219;
assign w7116 = (w6130 & ~w6287) | (w6130 & w16364) | (~w6287 & w16364);
assign w7117 = (w6174 & ~w6357) | (w6174 & w17619) | (~w6357 & w17619);
assign w7118 = ~w3683 & w7117;
assign w7119 = (~w6098 & ~w5470) | (~w6098 & w18034) | (~w5470 & w18034);
assign w7120 = ~w5224 & w6580;
assign w7121 = (w6143 & ~w6194) | (w6143 & w17156) | (~w6194 & w17156);
assign w7122 = w6134 & ~w6262;
assign w7123 = w6146 & ~w6381;
assign w7124 = (~w7119 & ~w6139) | (~w7119 & w16365) | (~w6139 & w16365);
assign w7125 = ~w6412 & w7124;
assign w7126 = ~w7116 & ~w7121;
assign w7127 = ~w7122 & w7126;
assign w7128 = ~w7115 & w7125;
assign w7129 = ~w7120 & ~w7123;
assign w7130 = w7128 & w7129;
assign w7131 = ~w7118 & w7127;
assign w7132 = w7130 & w7131;
assign w7133 = pi016 & w7132;
assign w7134 = ~w2723 & w6232;
assign w7135 = ~w6219 & w7134;
assign w7136 = ~w1137 & w6382;
assign w7137 = ~w3623 & w6174;
assign w7138 = (w7137 & ~w6357) | (w7137 & w17620) | (~w6357 & w17620);
assign w7139 = w2416 & w6159;
assign w7140 = (w7139 & ~w6257) | (w7139 & w16366) | (~w6257 & w16366);
assign w7141 = w4400 & w5632;
assign w7142 = (w7141 & ~w6287) | (w7141 & w16367) | (~w6287 & w16367);
assign w7143 = ~w7140 & ~w7142;
assign w7144 = ~w7138 & w7143;
assign w7145 = ~w7136 & w7144;
assign w7146 = (w5645 & ~w6194) | (w5645 & w18323) | (~w6194 & w18323);
assign w7147 = (w16368 & ~w6194) | (w16368 & w17157) | (~w6194 & w17157);
assign w7148 = (~w5857 & ~w5470) | (~w5857 & w18035) | (~w5470 & w18035);
assign w7149 = w6139 & w16369;
assign w7150 = ~w6426 & w7149;
assign w7151 = ~w7147 & w7150;
assign w7152 = w7150 & w17158;
assign w7153 = w7145 & w7152;
assign w7154 = w6963 & w6970;
assign w7155 = w4739 & w7154;
assign w7156 = w6695 & w7155;
assign w7157 = w7153 & w7156;
assign w7158 = pi018 & w7157;
assign w7159 = ~w6417 & ~w7114;
assign w7160 = ~w6694 & ~w7133;
assign w7161 = w7159 & w7160;
assign w7162 = ~w7158 & w7161;
assign w7163 = ~w6693 & w7162;
assign w7164 = (~w6392 & ~w7131) | (~w6392 & w17879) | (~w7131 & w17879);
assign w7165 = ~w6219 & w6232;
assign w7166 = (w7165 & ~w6557) | (w7165 & w16370) | (~w6557 & w16370);
assign w7167 = ~w2961 & w7166;
assign w7168 = w6934 & ~w7113;
assign w7169 = (w6380 & ~w6330) | (w6380 & w17621) | (~w6330 & w17621);
assign w7170 = ~w6650 & w7169;
assign w7171 = w6636 & w7170;
assign w7172 = w6649 & w7171;
assign w7173 = (w6382 & ~w6649) | (w6382 & w16371) | (~w6649 & w16371);
assign w7174 = w6382 & w18469;
assign w7175 = (w6580 & ~w6440) | (w6580 & w16372) | (~w6440 & w16372);
assign w7176 = ~w5253 & w7175;
assign w7177 = (w6561 & ~w6194) | (w6561 & w18037) | (~w6194 & w18037);
assign w7178 = ~w4854 & w6588;
assign w7179 = w6565 & w7178;
assign w7180 = w3404 & w7179;
assign w7181 = w7177 & w7180;
assign w7182 = w6585 & w7181;
assign w7183 = w6576 & w7182;
assign w7184 = (w7146 & ~w7182) | (w7146 & w17159) | (~w7182 & w17159);
assign w7185 = w628 & w7184;
assign w7186 = (~w6307 & ~w6684) | (~w6307 & w17160) | (~w6684 & w17160);
assign w7187 = ~w2134 & w6406;
assign w7188 = (w7187 & ~w6607) | (w7187 & w16373) | (~w6607 & w16373);
assign w7189 = w6389 & w7154;
assign w7190 = (w7189 & w6219) | (w7189 & w18038) | (w6219 & w18038);
assign w7191 = w7151 & w7190;
assign w7192 = w7145 & w7191;
assign w7193 = (w6963 & ~w7145) | (w6963 & w17622) | (~w7145 & w17622);
assign w7194 = ~w5799 & ~w6128;
assign w7195 = (w7194 & ~w6403) | (w7194 & w16374) | (~w6403 & w16374);
assign w7196 = (w7117 & ~w6485) | (w7117 & w17161) | (~w6485 & w17161);
assign w7197 = ~w3595 & w7196;
assign w7198 = (w6450 & ~w16345) | (w6450 & w17162) | (~w16345 & w17162);
assign w7199 = ~w4342 & w7198;
assign w7200 = w7089 & w7168;
assign w7201 = ~w7164 & w7200;
assign w7202 = ~w7186 & ~w7188;
assign w7203 = ~w7193 & ~w7195;
assign w7204 = w7202 & w7203;
assign w7205 = ~w7167 & w7201;
assign w7206 = ~w7174 & ~w7176;
assign w7207 = w7205 & w7206;
assign w7208 = ~w7185 & w7204;
assign w7209 = ~w7197 & ~w7199;
assign w7210 = w7208 & w7209;
assign w7211 = w7207 & w7210;
assign w7212 = pi017 & w7211;
assign w7213 = (w6451 & ~w16345) | (w6451 & w17163) | (~w16345 & w17163);
assign w7214 = (w6412 & ~w6461) | (w6412 & w17164) | (~w6461 & w17164);
assign w7215 = (w17159 & w17623) | (w17159 & w17624) | (w17623 & w17624);
assign w7216 = ~w7186 & w7214;
assign w7217 = ~w7213 & w7216;
assign w7218 = ~w7215 & w7217;
assign w7219 = (w6452 & ~w6485) | (w6452 & w17165) | (~w6485 & w17165);
assign w7220 = (w6455 & ~w6557) | (w6455 & w17625) | (~w6557 & w17625);
assign w7221 = ~w7219 & ~w7220;
assign w7222 = (w6406 & ~w6607) | (w6406 & w16375) | (~w6607 & w16375);
assign w7223 = w6406 & w18470;
assign w7224 = (w6454 & ~w6649) | (w6454 & w16376) | (~w6649 & w16376);
assign w7225 = (w6448 & ~w6440) | (w6448 & w16377) | (~w6440 & w16377);
assign w7226 = ~w7224 & ~w7225;
assign w7227 = ~w7223 & w7226;
assign w7228 = w7221 & w7227;
assign w7229 = w7218 & w7228;
assign w7230 = pi014 & w7229;
assign w7231 = pi183 & ~pi199;
assign w7232 = ~pi183 & pi199;
assign w7233 = pi184 & ~pi200;
assign w7234 = ~pi184 & pi200;
assign w7235 = pi185 & ~pi201;
assign w7236 = ~pi185 & pi201;
assign w7237 = ~pi186 & pi202;
assign w7238 = pi186 & ~pi202;
assign w7239 = pi187 & ~pi203;
assign w7240 = ~pi187 & pi203;
assign w7241 = ~pi188 & pi204;
assign w7242 = pi188 & ~pi204;
assign w7243 = pi189 & ~pi205;
assign w7244 = ~pi189 & pi205;
assign w7245 = pi190 & ~pi206;
assign w7246 = ~w7244 & w7245;
assign w7247 = ~w7242 & ~w7243;
assign w7248 = ~w7246 & w7247;
assign w7249 = ~w7240 & ~w7241;
assign w7250 = ~w7248 & w7249;
assign w7251 = ~w7238 & ~w7239;
assign w7252 = ~w7250 & w7251;
assign w7253 = ~w7236 & ~w7237;
assign w7254 = ~w7252 & w7253;
assign w7255 = ~w7235 & ~w7254;
assign w7256 = ~w7234 & ~w7255;
assign w7257 = ~w7233 & ~w7256;
assign w7258 = ~w7232 & ~w7257;
assign w7259 = ~w7231 & ~w7258;
assign w7260 = pi183 & ~pi223;
assign w7261 = ~pi183 & pi223;
assign w7262 = pi184 & ~pi224;
assign w7263 = ~pi184 & pi224;
assign w7264 = pi185 & ~pi225;
assign w7265 = ~pi185 & pi225;
assign w7266 = pi186 & ~pi226;
assign w7267 = ~pi186 & pi226;
assign w7268 = pi187 & ~pi227;
assign w7269 = ~pi187 & pi227;
assign w7270 = ~pi188 & pi228;
assign w7271 = pi189 & ~pi229;
assign w7272 = ~pi189 & pi229;
assign w7273 = pi190 & ~pi230;
assign w7274 = ~w7272 & w7273;
assign w7275 = ~w7271 & ~w7274;
assign w7276 = ~w7270 & ~w7275;
assign w7277 = pi188 & ~pi228;
assign w7278 = ~w7276 & ~w7277;
assign w7279 = ~w7269 & ~w7278;
assign w7280 = ~w7268 & ~w7279;
assign w7281 = ~w7267 & ~w7280;
assign w7282 = ~w7266 & ~w7281;
assign w7283 = ~w7265 & ~w7282;
assign w7284 = ~w7264 & ~w7283;
assign w7285 = ~w7263 & ~w7284;
assign w7286 = ~w7262 & ~w7285;
assign w7287 = ~w7261 & ~w7286;
assign w7288 = ~w7260 & ~w7287;
assign w7289 = pi183 & ~pi215;
assign w7290 = ~pi183 & pi215;
assign w7291 = pi184 & ~pi216;
assign w7292 = ~pi184 & pi216;
assign w7293 = pi185 & ~pi217;
assign w7294 = ~pi186 & pi218;
assign w7295 = ~pi185 & pi217;
assign w7296 = pi186 & ~pi218;
assign w7297 = ~pi187 & pi219;
assign w7298 = pi187 & ~pi219;
assign w7299 = ~pi188 & pi220;
assign w7300 = pi188 & ~pi220;
assign w7301 = ~pi189 & pi221;
assign w7302 = pi189 & ~pi221;
assign w7303 = pi190 & ~pi222;
assign w7304 = ~w7302 & ~w7303;
assign w7305 = ~w7301 & ~w7304;
assign w7306 = ~w7300 & ~w7305;
assign w7307 = ~w7299 & ~w7306;
assign w7308 = ~w7298 & ~w7307;
assign w7309 = ~w7297 & ~w7308;
assign w7310 = ~w7296 & ~w7309;
assign w7311 = ~w7294 & ~w7295;
assign w7312 = ~w7310 & w7311;
assign w7313 = ~w7293 & ~w7312;
assign w7314 = ~w7292 & ~w7313;
assign w7315 = ~w7291 & ~w7314;
assign w7316 = ~w7290 & ~w7315;
assign w7317 = ~w7289 & ~w7316;
assign w7318 = w7288 & w7317;
assign w7319 = pi183 & ~pi207;
assign w7320 = ~pi183 & pi207;
assign w7321 = pi184 & ~pi208;
assign w7322 = ~pi184 & pi208;
assign w7323 = pi185 & ~pi209;
assign w7324 = ~pi185 & pi209;
assign w7325 = pi186 & ~pi210;
assign w7326 = ~pi186 & pi210;
assign w7327 = pi187 & ~pi211;
assign w7328 = ~pi187 & pi211;
assign w7329 = ~pi188 & pi212;
assign w7330 = pi189 & ~pi213;
assign w7331 = ~pi189 & pi213;
assign w7332 = pi190 & ~pi214;
assign w7333 = ~w7331 & w7332;
assign w7334 = ~w7330 & ~w7333;
assign w7335 = ~w7329 & ~w7334;
assign w7336 = pi188 & ~pi212;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = ~w7328 & ~w7337;
assign w7339 = ~w7327 & ~w7338;
assign w7340 = ~w7326 & ~w7339;
assign w7341 = ~w7325 & ~w7340;
assign w7342 = ~w7324 & ~w7341;
assign w7343 = ~w7323 & ~w7342;
assign w7344 = ~w7322 & ~w7343;
assign w7345 = ~w7321 & ~w7344;
assign w7346 = ~w7320 & ~w7345;
assign w7347 = ~w7319 & ~w7346;
assign w7348 = w7259 & w7347;
assign w7349 = w7318 & w7348;
assign w7350 = ~pi183 & pi239;
assign w7351 = pi183 & ~pi239;
assign w7352 = ~pi184 & pi240;
assign w7353 = pi184 & ~pi240;
assign w7354 = ~pi185 & pi241;
assign w7355 = pi186 & ~pi242;
assign w7356 = pi185 & ~pi241;
assign w7357 = ~pi186 & pi242;
assign w7358 = pi187 & ~pi243;
assign w7359 = ~pi187 & pi243;
assign w7360 = pi189 & ~pi245;
assign w7361 = ~pi189 & pi245;
assign w7362 = pi190 & ~pi246;
assign w7363 = ~w7361 & w7362;
assign w7364 = ~w7360 & ~w7363;
assign w7365 = pi244 & w7364;
assign w7366 = pi188 & ~w7365;
assign w7367 = ~pi244 & ~w7364;
assign w7368 = ~w7366 & ~w7367;
assign w7369 = ~w7359 & ~w7368;
assign w7370 = ~w7358 & ~w7369;
assign w7371 = ~w7357 & ~w7370;
assign w7372 = ~w7355 & ~w7356;
assign w7373 = ~w7371 & w7372;
assign w7374 = ~w7354 & ~w7373;
assign w7375 = ~w7353 & ~w7374;
assign w7376 = ~w7352 & ~w7375;
assign w7377 = ~w7351 & ~w7376;
assign w7378 = ~w7350 & ~w7377;
assign w7379 = ~pi183 & pi255;
assign w7380 = pi183 & ~pi255;
assign w7381 = ~pi184 & pi256;
assign w7382 = pi184 & ~pi256;
assign w7383 = ~pi185 & pi257;
assign w7384 = pi185 & ~pi257;
assign w7385 = pi186 & ~pi258;
assign w7386 = ~pi186 & pi258;
assign w7387 = ~pi187 & pi259;
assign w7388 = pi189 & ~pi261;
assign w7389 = ~pi189 & pi261;
assign w7390 = pi190 & ~pi262;
assign w7391 = ~w7389 & w7390;
assign w7392 = ~w7388 & ~w7391;
assign w7393 = ~pi260 & ~w7392;
assign w7394 = pi187 & ~pi259;
assign w7395 = pi260 & w7392;
assign w7396 = pi188 & ~w7395;
assign w7397 = ~w7393 & ~w7394;
assign w7398 = ~w7396 & w7397;
assign w7399 = ~w7386 & ~w7387;
assign w7400 = ~w7398 & w7399;
assign w7401 = ~w7384 & ~w7385;
assign w7402 = ~w7400 & w7401;
assign w7403 = ~w7383 & ~w7402;
assign w7404 = ~w7382 & ~w7403;
assign w7405 = ~w7381 & ~w7404;
assign w7406 = ~w7380 & ~w7405;
assign w7407 = ~w7379 & ~w7406;
assign w7408 = pi183 & ~pi263;
assign w7409 = ~pi183 & pi263;
assign w7410 = pi184 & ~pi264;
assign w7411 = ~pi184 & pi264;
assign w7412 = pi185 & ~pi265;
assign w7413 = ~pi185 & pi265;
assign w7414 = pi186 & ~pi266;
assign w7415 = ~pi186 & pi266;
assign w7416 = pi187 & ~pi267;
assign w7417 = ~pi187 & pi267;
assign w7418 = ~pi188 & pi268;
assign w7419 = pi189 & ~pi269;
assign w7420 = ~pi189 & pi269;
assign w7421 = pi190 & ~pi270;
assign w7422 = ~w7420 & w7421;
assign w7423 = ~w7419 & ~w7422;
assign w7424 = ~w7418 & ~w7423;
assign w7425 = pi188 & ~pi268;
assign w7426 = ~w7424 & ~w7425;
assign w7427 = ~w7417 & ~w7426;
assign w7428 = ~w7416 & ~w7427;
assign w7429 = ~w7415 & ~w7428;
assign w7430 = ~w7414 & ~w7429;
assign w7431 = ~w7413 & ~w7430;
assign w7432 = ~w7412 & ~w7431;
assign w7433 = ~w7411 & ~w7432;
assign w7434 = ~w7410 & ~w7433;
assign w7435 = ~w7409 & ~w7434;
assign w7436 = ~w7408 & ~w7435;
assign w7437 = pi183 & ~pi271;
assign w7438 = ~pi183 & pi271;
assign w7439 = pi184 & ~pi272;
assign w7440 = ~pi184 & pi272;
assign w7441 = pi185 & ~pi273;
assign w7442 = ~pi185 & pi273;
assign w7443 = ~pi186 & pi274;
assign w7444 = pi186 & ~pi274;
assign w7445 = pi187 & ~pi275;
assign w7446 = ~pi187 & pi275;
assign w7447 = ~pi188 & pi276;
assign w7448 = pi188 & ~pi276;
assign w7449 = pi189 & ~pi277;
assign w7450 = ~pi189 & pi277;
assign w7451 = pi190 & ~pi278;
assign w7452 = ~w7450 & w7451;
assign w7453 = ~w7448 & ~w7449;
assign w7454 = ~w7452 & w7453;
assign w7455 = ~w7446 & ~w7447;
assign w7456 = ~w7454 & w7455;
assign w7457 = ~w7444 & ~w7445;
assign w7458 = ~w7456 & w7457;
assign w7459 = ~w7442 & ~w7443;
assign w7460 = ~w7458 & w7459;
assign w7461 = ~w7441 & ~w7460;
assign w7462 = ~w7440 & ~w7461;
assign w7463 = ~w7439 & ~w7462;
assign w7464 = ~w7438 & ~w7463;
assign w7465 = ~w7437 & ~w7464;
assign w7466 = w7436 & w7465;
assign w7467 = pi183 & ~pi247;
assign w7468 = ~pi183 & pi247;
assign w7469 = pi184 & ~pi248;
assign w7470 = ~pi184 & pi248;
assign w7471 = pi185 & ~pi249;
assign w7472 = ~pi186 & pi250;
assign w7473 = ~pi185 & pi249;
assign w7474 = pi186 & ~pi250;
assign w7475 = ~pi187 & pi251;
assign w7476 = pi187 & ~pi251;
assign w7477 = ~pi188 & pi252;
assign w7478 = pi188 & ~pi252;
assign w7479 = ~pi189 & pi253;
assign w7480 = pi189 & ~pi253;
assign w7481 = pi190 & ~pi254;
assign w7482 = ~w7480 & ~w7481;
assign w7483 = ~w7479 & ~w7482;
assign w7484 = ~w7478 & ~w7483;
assign w7485 = ~w7477 & ~w7484;
assign w7486 = ~w7476 & ~w7485;
assign w7487 = ~w7475 & ~w7486;
assign w7488 = ~w7474 & ~w7487;
assign w7489 = ~w7472 & ~w7473;
assign w7490 = ~w7488 & w7489;
assign w7491 = ~w7471 & ~w7490;
assign w7492 = ~w7470 & ~w7491;
assign w7493 = ~w7469 & ~w7492;
assign w7494 = ~w7468 & ~w7493;
assign w7495 = ~w7467 & ~w7494;
assign w7496 = ~w7407 & w7495;
assign w7497 = w7466 & w7496;
assign w7498 = pi183 & ~pi231;
assign w7499 = ~pi183 & pi231;
assign w7500 = pi184 & ~pi232;
assign w7501 = ~pi184 & pi232;
assign w7502 = pi185 & ~pi233;
assign w7503 = ~pi185 & pi233;
assign w7504 = pi186 & ~pi234;
assign w7505 = ~pi186 & pi234;
assign w7506 = pi187 & ~pi235;
assign w7507 = ~pi187 & pi235;
assign w7508 = ~pi188 & pi236;
assign w7509 = pi189 & ~pi237;
assign w7510 = ~pi189 & pi237;
assign w7511 = pi190 & ~pi238;
assign w7512 = ~w7510 & w7511;
assign w7513 = ~w7509 & ~w7512;
assign w7514 = ~w7508 & ~w7513;
assign w7515 = pi188 & ~pi236;
assign w7516 = ~w7514 & ~w7515;
assign w7517 = ~w7507 & ~w7516;
assign w7518 = ~w7506 & ~w7517;
assign w7519 = ~w7505 & ~w7518;
assign w7520 = ~w7504 & ~w7519;
assign w7521 = ~w7503 & ~w7520;
assign w7522 = ~w7502 & ~w7521;
assign w7523 = ~w7501 & ~w7522;
assign w7524 = ~w7500 & ~w7523;
assign w7525 = ~w7499 & ~w7524;
assign w7526 = ~w7498 & ~w7525;
assign w7527 = ~w7378 & w7526;
assign w7528 = w7497 & w7527;
assign w7529 = w4724 & w7107;
assign w7530 = ~w823 & w7529;
assign w7531 = ~pi183 & ~w6935;
assign w7532 = w4726 & w7531;
assign w7533 = ~w7530 & ~w7532;
assign w7534 = ~w693 & w4730;
assign w7535 = w2597 & w7534;
assign w7536 = w6970 & w7535;
assign w7537 = pi183 & ~pi191;
assign w7538 = ~pi183 & pi191;
assign w7539 = pi184 & ~pi192;
assign w7540 = ~pi184 & pi192;
assign w7541 = pi185 & ~pi193;
assign w7542 = ~pi185 & pi193;
assign w7543 = ~pi186 & pi194;
assign w7544 = pi186 & ~pi194;
assign w7545 = pi187 & ~pi195;
assign w7546 = ~pi187 & pi195;
assign w7547 = ~pi188 & pi196;
assign w7548 = pi188 & ~pi196;
assign w7549 = pi189 & ~pi197;
assign w7550 = ~pi189 & pi197;
assign w7551 = pi190 & ~pi198;
assign w7552 = ~w7550 & w7551;
assign w7553 = ~w7548 & ~w7549;
assign w7554 = ~w7552 & w7553;
assign w7555 = ~w7546 & ~w7547;
assign w7556 = ~w7554 & w7555;
assign w7557 = ~w7544 & ~w7545;
assign w7558 = ~w7556 & w7557;
assign w7559 = ~w7542 & ~w7543;
assign w7560 = ~w7558 & w7559;
assign w7561 = ~w7541 & ~w7560;
assign w7562 = ~w7540 & ~w7561;
assign w7563 = ~w7539 & ~w7562;
assign w7564 = ~w7538 & ~w7563;
assign w7565 = ~w7537 & ~w7564;
assign w7566 = ~w6097 & ~w6962;
assign w7567 = ~w2040 & ~w7533;
assign w7568 = w7536 & w7567;
assign w7569 = w821 & w7568;
assign w7570 = w2546 & ~w3223;
assign w7571 = ~w5827 & ~w7086;
assign w7572 = w7570 & w7571;
assign w7573 = ~w1668 & w7569;
assign w7574 = w4551 & w4717;
assign w7575 = w7566 & w7574;
assign w7576 = w7572 & w7573;
assign w7577 = w6100 & w7576;
assign w7578 = w7565 & w7575;
assign w7579 = w7577 & w7578;
assign w7580 = w6106 & w7579;
assign w7581 = ~w5192 & w7580;
assign w7582 = w7349 & w7581;
assign w7583 = w7528 & w7582;
assign w7584 = w7145 & w17626;
assign w7585 = w3949 & w7584;
assign w7586 = pi019 & w7585;
assign w7587 = (w7118 & ~w6485) | (w7118 & w18324) | (~w6485 & w18324);
assign w7588 = (w7116 & ~w16345) | (w7116 & w18040) | (~w16345 & w18040);
assign w7589 = (w7122 & ~w6607) | (w7122 & w16378) | (~w6607 & w16378);
assign w7590 = (w7120 & ~w6440) | (w7120 & w16379) | (~w6440 & w16379);
assign w7591 = w691 & w7184;
assign w7592 = (w7115 & ~w6557) | (w7115 & w16380) | (~w6557 & w16380);
assign w7593 = (w7119 & ~w6403) | (w7119 & w16381) | (~w6403 & w16381);
assign w7594 = w6382 & w18471;
assign w7595 = w7164 & ~w7214;
assign w7596 = ~w7589 & ~w7590;
assign w7597 = ~w7592 & ~w7593;
assign w7598 = w7596 & w7597;
assign w7599 = ~w7587 & w7595;
assign w7600 = ~w7588 & ~w7594;
assign w7601 = w7599 & w7600;
assign w7602 = ~w7591 & w7598;
assign w7603 = w7601 & w7602;
assign w7604 = pi016 & w7603;
assign w7605 = w6406 & w18472;
assign w7606 = (~w6963 & ~w6149) | (~w6963 & w18043) | (~w6149 & w18043);
assign w7607 = (w7148 & ~w6403) | (w7148 & w16382) | (~w6403 & w16382);
assign w7608 = (w16383 & w7135) | (w16383 & w18044) | (w7135 & w18044);
assign w7609 = (w7136 & ~w6649) | (w7136 & w16384) | (~w6649 & w16384);
assign w7610 = (w7142 & ~w16345) | (w7142 & w17166) | (~w16345 & w17166);
assign w7611 = (~w6440 & w17627) | (~w6440 & w17628) | (w17627 & w17628);
assign w7612 = (w7138 & ~w6485) | (w7138 & w17167) | (~w6485 & w17167);
assign w7613 = (w7147 & ~w7182) | (w7147 & w17168) | (~w7182 & w17168);
assign w7614 = ~w5431 & ~w7606;
assign w7615 = (w7614 & ~w7145) | (w7614 & w17629) | (~w7145 & w17629);
assign w7616 = ~w7164 & w7615;
assign w7617 = ~w7607 & ~w7609;
assign w7618 = w7616 & w7617;
assign w7619 = ~w7605 & ~w7608;
assign w7620 = ~w7610 & ~w7611;
assign w7621 = ~w7612 & ~w7613;
assign w7622 = w7620 & w7621;
assign w7623 = w7618 & w7619;
assign w7624 = w7622 & w7623;
assign w7625 = pi018 & w7624;
assign w7626 = (w17159 & w17630) | (w17159 & w17631) | (w17630 & w17631);
assign w7627 = w7189 & ~w7565;
assign w7628 = ~w7626 & w7627;
assign w7629 = w6450 & w18473;
assign w7630 = ~w6999 & ~w7113;
assign w7631 = ~w5282 & w6580;
assign w7632 = (w7631 & ~w6440) | (w7631 & w16385) | (~w6440 & w16385);
assign w7633 = w5769 & ~w6128;
assign w7634 = (w7633 & ~w6403) | (w7633 & w17633) | (~w6403 & w17633);
assign w7635 = w3565 & w7117;
assign w7636 = (w7635 & ~w6485) | (w7635 & w17169) | (~w6485 & w17169);
assign w7637 = (w16371 & w18045) | (w16371 & w18046) | (w18045 & w18046);
assign w7638 = (w16370 & w17170) | (w16370 & w17171) | (w17170 & w17171);
assign w7639 = (w16375 & w18047) | (w16375 & w18048) | (w18047 & w18048);
assign w7640 = w7145 & w17172;
assign w7641 = ~w7632 & w7640;
assign w7642 = ~w7634 & w7641;
assign w7643 = ~w7636 & ~w7637;
assign w7644 = ~w7638 & ~w7639;
assign w7645 = w7643 & w7644;
assign w7646 = ~w7629 & w7642;
assign w7647 = w7645 & w7646;
assign w7648 = w7646 & w18049;
assign w7649 = pi020 & w7648;
assign w7650 = (w6395 & ~w16345) | (w6395 & w17173) | (~w16345 & w17173);
assign w7651 = (w6397 & ~w6440) | (w6397 & w17634) | (~w6440 & w17634);
assign w7652 = w6399 & ~w7183;
assign w7653 = (w6393 & ~w7131) | (w6393 & w18050) | (~w7131 & w18050);
assign w7654 = (w6410 & ~w6557) | (w6410 & w17635) | (~w6557 & w17635);
assign w7655 = w5799 & ~w7113;
assign w7656 = (~w5828 & ~w6403) | (~w5828 & w17636) | (~w6403 & w17636);
assign w7657 = (~w17164 & w17637) | (~w17164 & w17638) | (w17637 & w17638);
assign w7658 = ~w7651 & ~w7653;
assign w7659 = ~w7654 & w7656;
assign w7660 = w7658 & w7659;
assign w7661 = ~w7650 & w7657;
assign w7662 = ~w7652 & w7661;
assign w7663 = w7660 & w7662;
assign w7664 = (w6383 & ~w6649) | (w6383 & w16386) | (~w6649 & w16386);
assign w7665 = (w6407 & ~w6607) | (w6407 & w16387) | (~w6607 & w16387);
assign w7666 = (w5857 & ~w7145) | (w5857 & w17639) | (~w7145 & w17639);
assign w7667 = w6405 & ~w6494;
assign w7668 = ~w7664 & ~w7665;
assign w7669 = ~w7666 & w7668;
assign w7670 = ~w7667 & w7669;
assign w7671 = w7663 & w7670;
assign w7672 = w5770 & w7671;
assign w7673 = w6376 & w7672;
assign w7674 = (w6423 & ~w6461) | (w6423 & w17174) | (~w6461 & w17174);
assign w7675 = (w6421 & ~w6649) | (w6421 & w16388) | (~w6649 & w16388);
assign w7676 = (w6422 & ~w6557) | (w6422 & w16389) | (~w6557 & w16389);
assign w7677 = ~w3714 & w7196;
assign w7678 = w5253 & ~w7113;
assign w7679 = w5341 & ~w7192;
assign w7680 = (w6419 & ~w6403) | (w6419 & w16390) | (~w6403 & w16390);
assign w7681 = w6418 & ~w7183;
assign w7682 = (w6429 & ~w6607) | (w6429 & w16391) | (~w6607 & w16391);
assign w7683 = (w6424 & ~w7131) | (w6424 & w18051) | (~w7131 & w18051);
assign w7684 = (w6428 & ~w16345) | (w6428 & w18325) | (~w16345 & w18325);
assign w7685 = w6420 & ~w7678;
assign w7686 = ~w7186 & w7685;
assign w7687 = w7632 & ~w7674;
assign w7688 = ~w7675 & ~w7676;
assign w7689 = ~w7679 & ~w7680;
assign w7690 = ~w7682 & ~w7683;
assign w7691 = w7689 & w7690;
assign w7692 = w7687 & w7688;
assign w7693 = ~w7681 & w7686;
assign w7694 = ~w7684 & w7693;
assign w7695 = w7691 & w16392;
assign w7696 = w7694 & w7695;
assign w7697 = ~pi013 & w7696;
assign w7698 = ~w5431 & w6375;
assign w7699 = w5770 & w7698;
assign w7700 = w7669 & w17640;
assign w7701 = w7663 & w7700;
assign w7702 = ~w7229 & ~w7701;
assign w7703 = w4342 & ~w7113;
assign w7704 = w6496 & ~w6685;
assign w7705 = (w6500 & ~w16347) | (w6500 & w17175) | (~w16347 & w17175);
assign w7706 = ~w1292 & w7173;
assign w7707 = w4371 & ~w7703;
assign w7708 = w7707 & w18474;
assign w7709 = ~w7704 & ~w7705;
assign w7710 = w7708 & w7709;
assign w7711 = ~w7706 & w7710;
assign w7712 = w4669 & w6289;
assign w7713 = (w6503 & ~w7131) | (w6503 & w17880) | (~w7131 & w17880);
assign w7714 = (w6502 & ~w6607) | (w6502 & w16393) | (~w6607 & w16393);
assign w7715 = w6505 & ~w7183;
assign w7716 = (w6497 & ~w6485) | (w6497 & w18052) | (~w6485 & w18052);
assign w7717 = (w16370 & w18053) | (w16370 & w18054) | (w18053 & w18054);
assign w7718 = w4163 & w7214;
assign w7719 = (w6506 & ~w6403) | (w6506 & w18055) | (~w6403 & w18055);
assign w7720 = w4134 & w7175;
assign w7721 = ~w7713 & ~w7714;
assign w7722 = ~w7719 & w7721;
assign w7723 = ~w7715 & ~w7716;
assign w7724 = ~w7717 & ~w7718;
assign w7725 = ~w7720 & w7724;
assign w7726 = w7722 & w7723;
assign w7727 = w7725 & w7726;
assign w7728 = ~w6523 & w7712;
assign w7729 = w7711 & w7728;
assign w7730 = w7727 & w7729;
assign w7731 = ~w4551 & w7730;
assign w7732 = w4461 & w6276;
assign w7733 = ~w6294 & w7732;
assign w7734 = ~pi011 & ~w4580;
assign w7735 = w7733 & w7734;
assign w7736 = w7731 & w7735;
assign w7737 = (w6676 & ~w16345) | (w6676 & w17176) | (~w16345 & w17176);
assign w7738 = (w16370 & w17177) | (w16370 & w17178) | (w17177 & w17178);
assign w7739 = ~w7737 & ~w7738;
assign w7740 = w2229 & w7222;
assign w7741 = (w6673 & ~w7182) | (w6673 & w17179) | (~w7182 & w17179);
assign w7742 = (w6678 & ~w6485) | (w6678 & w17180) | (~w6485 & w17180);
assign w7743 = (w6677 & ~w6649) | (w6677 & w17642) | (~w6649 & w17642);
assign w7744 = ~w6685 & ~w7705;
assign w7745 = ~w7743 & w7744;
assign w7746 = ~w7741 & ~w7742;
assign w7747 = w7745 & w7746;
assign w7748 = (~w5431 & w17643) | (~w5431 & ~w7222) | (w17643 & ~w7222);
assign w7749 = w7739 & w7748;
assign w7750 = w7747 & w7749;
assign w7751 = ~w6307 & w7750;
assign w7752 = ~w6517 & w6522;
assign w7753 = w7710 & w18326;
assign w7754 = w7727 & w7753;
assign w7755 = ~w1417 & w7173;
assign w7756 = (w6473 & ~w6440) | (w6473 & w16394) | (~w6440 & w16394);
assign w7757 = ~w6466 & ~w6533;
assign w7758 = w6342 & w7186;
assign w7759 = ~w7757 & ~w7758;
assign w7760 = (w6476 & ~w6403) | (w6476 & w16395) | (~w6403 & w16395);
assign w7761 = (w6469 & ~w6557) | (w6469 & w16396) | (~w6557 & w16396);
assign w7762 = (w6488 & ~w7131) | (w6488 & w17881) | (~w7131 & w17881);
assign w7763 = (w6489 & ~w6607) | (w6489 & w16397) | (~w6607 & w16397);
assign w7764 = ~w6462 & w6487;
assign w7765 = (w3623 & ~w7145) | (w3623 & w17644) | (~w7145 & w17644);
assign w7766 = w3595 & ~w7113;
assign w7767 = (w6440 & w18056) | (w6440 & w18057) | (w18056 & w18057);
assign w7768 = ~w7760 & ~w7761;
assign w7769 = ~w7762 & ~w7763;
assign w7770 = ~w7764 & ~w7765;
assign w7771 = w7769 & w7770;
assign w7772 = w7767 & w7768;
assign w7773 = ~w7755 & w7772;
assign w7774 = w7759 & w7771;
assign w7775 = w7773 & w7774;
assign w7776 = ~w278 & w7184;
assign w7777 = w4009 & w7198;
assign w7778 = ~w7776 & ~w7777;
assign w7779 = w3536 & ~w3949;
assign w7780 = w3920 & w7779;
assign w7781 = w7636 & w7780;
assign w7782 = w7778 & w7781;
assign w7783 = w7775 & w7782;
assign w7784 = ~pi009 & w7783;
assign w7785 = (w17159 & w17645) | (w17159 & w17646) | (w17645 & w17646);
assign w7786 = w6382 & w18475;
assign w7787 = (w6524 & ~w6557) | (w6524 & w16398) | (~w6557 & w16398);
assign w7788 = (w6528 & ~w6607) | (w6528 & w16399) | (~w6607 & w16399);
assign w7789 = (w6527 & ~w6485) | (w6527 & w17181) | (~w6485 & w17181);
assign w7790 = ~w6464 & w7705;
assign w7791 = ~w7787 & ~w7788;
assign w7792 = w7790 & w7791;
assign w7793 = ~w7786 & ~w7789;
assign w7794 = w7792 & w7793;
assign w7795 = w7792 & w17182;
assign w7796 = (w6544 & ~w16347) | (w6544 & w17183) | (~w16347 & w17183);
assign w7797 = w3258 & w6225;
assign w7798 = ~w7796 & ~w7797;
assign w7799 = (w6535 & ~w6649) | (w6535 & w16400) | (~w6649 & w16400);
assign w7800 = ~w6494 & w6546;
assign w7801 = (w6545 & ~w6403) | (w6545 & w16401) | (~w6403 & w16401);
assign w7802 = ~w7799 & ~w7801;
assign w7803 = w7798 & w7802;
assign w7804 = ~w7800 & w7803;
assign w7805 = ~w342 & w7184;
assign w7806 = w5525 & w7165;
assign w7807 = (w16402 & ~w7131) | (w16402 & w17882) | (~w7131 & w17882);
assign w7808 = (~w6440 & w17647) | (~w6440 & w17648) | (w17647 & w17648);
assign w7809 = (w6543 & ~w6607) | (w6543 & w17649) | (~w6607 & w17649);
assign w7810 = (w17164 & w17650) | (w17164 & w17651) | (w17650 & w17651);
assign w7811 = (w2723 & ~w7145) | (w2723 & w17652) | (~w7145 & w17652);
assign w7812 = (w6537 & ~w16345) | (w6537 & w17184) | (~w16345 & w17184);
assign w7813 = (w2961 & ~w6149) | (w2961 & w18058) | (~w6149 & w18058);
assign w7814 = w6548 & ~w6685;
assign w7815 = w6200 & ~w7813;
assign w7816 = (w7815 & ~w6557) | (w7815 & w17653) | (~w6557 & w17653);
assign w7817 = ~w7809 & w7816;
assign w7818 = ~w7811 & ~w7814;
assign w7819 = w7817 & w7818;
assign w7820 = ~w7807 & ~w7808;
assign w7821 = ~w7810 & ~w7812;
assign w7822 = w7820 & w7821;
assign w7823 = w7819 & w7822;
assign w7824 = w5526 & w7806;
assign w7825 = ~w7805 & w7824;
assign w7826 = w7804 & w7825;
assign w7827 = w7823 & w7826;
assign w7828 = pi007 & w7827;
assign w7829 = w2134 & ~w7113;
assign w7830 = w2322 & ~w7829;
assign w7831 = ~w6533 & w6596;
assign w7832 = (~w4797 & w6533) | (~w4797 & w18059) | (w6533 & w18059);
assign w7833 = (w6611 & ~w6403) | (w6611 & w16403) | (~w6403 & w16403);
assign w7834 = (w6601 & ~w6684) | (w6601 & w17185) | (~w6684 & w17185);
assign w7835 = ~w2416 & ~w7192;
assign w7836 = ~w7833 & ~w7834;
assign w7837 = ~w7835 & w7836;
assign w7838 = w7832 & w7837;
assign w7839 = ~w6628 & w6660;
assign w7840 = (w6608 & ~w6649) | (w6608 & w16404) | (~w6649 & w16404);
assign w7841 = (w6597 & ~w6440) | (w6597 & w16405) | (~w6440 & w16405);
assign w7842 = (w6599 & ~w7131) | (w6599 & w18060) | (~w7131 & w18060);
assign w7843 = (w16383 & w17186) | (w16383 & w17187) | (w17186 & w17187);
assign w7844 = (w17164 & w17654) | (w17164 & w17655) | (w17654 & w17655);
assign w7845 = (w6594 & ~w6485) | (w6594 & w17188) | (~w6485 & w17188);
assign w7846 = (w6598 & ~w16345) | (w6598 & w17189) | (~w16345 & w17189);
assign w7847 = w6609 & ~w7183;
assign w7848 = ~w7840 & ~w7841;
assign w7849 = ~w7842 & w7848;
assign w7850 = ~w7843 & ~w7844;
assign w7851 = ~w7845 & ~w7846;
assign w7852 = ~w7847 & w7851;
assign w7853 = w7849 & w7850;
assign w7854 = w7852 & w7853;
assign w7855 = w7830 & w7839;
assign w7856 = w7838 & w7855;
assign w7857 = w7854 & w7856;
assign w7858 = w6622 & w7857;
assign w7859 = w6664 & w7858;
assign w7860 = ~w628 & ~w7113;
assign w7861 = (w6560 & ~w6403) | (w6560 & w16406) | (~w6403 & w16406);
assign w7862 = w6571 & ~w6685;
assign w7863 = ~w6462 & w6572;
assign w7864 = (w6570 & ~w6649) | (w6570 & w16407) | (~w6649 & w16407);
assign w7865 = (w659 & ~w7145) | (w659 & w17656) | (~w7145 & w17656);
assign w7866 = (w6579 & ~w7131) | (w6579 & w17883) | (~w7131 & w17883);
assign w7867 = (w6578 & ~w6607) | (w6578 & w16408) | (~w6607 & w16408);
assign w7868 = (w6581 & ~w6440) | (w6581 & w16409) | (~w6440 & w16409);
assign w7869 = (w6568 & ~w6557) | (w6568 & w16410) | (~w6557 & w16410);
assign w7870 = (w6577 & ~w16345) | (w6577 & w17190) | (~w16345 & w17190);
assign w7871 = (w6569 & ~w6485) | (w6569 & w17191) | (~w6485 & w17191);
assign w7872 = (w6567 & ~w16347) | (w6567 & w17192) | (~w16347 & w17192);
assign w7873 = ~w6180 & ~w7872;
assign w7874 = ~w7183 & ~w7861;
assign w7875 = ~w7862 & ~w7863;
assign w7876 = ~w7864 & ~w7865;
assign w7877 = ~w7866 & ~w7867;
assign w7878 = ~w7868 & ~w7869;
assign w7879 = w7877 & w7878;
assign w7880 = w7875 & w7876;
assign w7881 = ~w7870 & w7874;
assign w7882 = ~w7871 & w7873;
assign w7883 = w7881 & w7882;
assign w7884 = w7879 & w7880;
assign w7885 = w7883 & w7884;
assign w7886 = w6588 & ~w7860;
assign w7887 = w7885 & w7886;
assign w7888 = ~w3337 & w6564;
assign w7889 = pi001 & w596;
assign w7890 = w7888 & w7889;
assign w7891 = w533 & ~w3346;
assign w7892 = w6562 & w7891;
assign w7893 = w220 & w7890;
assign w7894 = w7892 & w7893;
assign w7895 = w7887 & w7894;
assign w7896 = w6625 & w7830;
assign w7897 = ~w6628 & w7896;
assign w7898 = w7837 & w17193;
assign w7899 = w7854 & w7898;
assign w7900 = w6333 & w6630;
assign w7901 = ~w7172 & w7900;
assign w7902 = (w6637 & ~w6485) | (w6637 & w17194) | (~w6485 & w17194);
assign w7903 = (w6632 & ~w7182) | (w6632 & w17195) | (~w7182 & w17195);
assign w7904 = (w6643 & ~w6461) | (w6643 & w17196) | (~w6461 & w17196);
assign w7905 = (w6650 & ~w6557) | (w6650 & w17657) | (~w6557 & w17657);
assign w7906 = (w1073 & ~w6149) | (w1073 & w18328) | (~w6149 & w18328);
assign w7907 = (w6641 & ~w6607) | (w6641 & w17658) | (~w6607 & w17658);
assign w7908 = (w1137 & ~w7145) | (w1137 & w17659) | (~w7145 & w17659);
assign w7909 = (w6631 & ~w6403) | (w6631 & w17660) | (~w6403 & w17660);
assign w7910 = (w6633 & ~w7131) | (w6633 & w18061) | (~w7131 & w18061);
assign w7911 = ~w1168 & ~w7906;
assign w7912 = (~w17196 & w17661) | (~w17196 & w17662) | (w17661 & w17662);
assign w7913 = ~w7905 & ~w7907;
assign w7914 = ~w7908 & ~w7909;
assign w7915 = w7913 & w7914;
assign w7916 = ~w7902 & w7912;
assign w7917 = ~w7903 & ~w7910;
assign w7918 = w7916 & w7917;
assign w7919 = w7915 & w7918;
assign w7920 = (w6640 & ~w16347) | (w6640 & w17197) | (~w16347 & w17197);
assign w7921 = w6318 & ~w7920;
assign w7922 = (w6639 & ~w6440) | (w6639 & w16411) | (~w6440 & w16411);
assign w7923 = w6638 & ~w6685;
assign w7924 = (w6642 & ~w16345) | (w6642 & w17198) | (~w16345 & w17198);
assign w7925 = (w6440 & w17663) | (w6440 & w17664) | (w17663 & w17664);
assign w7926 = ~w7923 & w7925;
assign w7927 = w7921 & ~w7924;
assign w7928 = w7926 & w7927;
assign w7929 = w7901 & w7928;
assign w7930 = w7919 & w7929;
assign w7931 = w5565 & w7930;
assign w7932 = ~w7895 & ~w7899;
assign w7933 = ~w7931 & w7932;
assign w7934 = ~w7827 & ~w7859;
assign w7935 = ~w7933 & w7934;
assign w7936 = ~w7783 & ~w7828;
assign w7937 = ~w7935 & w7936;
assign w7938 = ~w7784 & ~w7795;
assign w7939 = ~w7937 & w7938;
assign w7940 = pi010 & w7795;
assign w7941 = ~w7754 & ~w7940;
assign w7942 = ~w7939 & w7941;
assign w7943 = ~w7736 & ~w7751;
assign w7944 = ~w7942 & w7943;
assign w7945 = pi012 & w7751;
assign w7946 = ~w7696 & ~w7945;
assign w7947 = ~w7944 & w7946;
assign w7948 = ~w7697 & w7702;
assign w7949 = ~w7947 & w7948;
assign w7950 = ~w7230 & ~w7586;
assign w7951 = ~w7604 & ~w7625;
assign w7952 = w7950 & w7951;
assign w7953 = ~w7212 & ~w7649;
assign w7954 = w7952 & w7953;
assign w7955 = ~w7673 & w7954;
assign w7956 = ~w7949 & w7955;
assign w7957 = (w7195 & ~w7663) | (w7195 & w17665) | (~w7663 & w17665);
assign w7958 = w6382 & w18476;
assign w7959 = w7927 & w17666;
assign w7960 = w7919 & w7959;
assign w7961 = (w7174 & ~w7919) | (w7174 & w17667) | (~w7919 & w17667);
assign w7962 = (w7197 & ~w7775) | (w7197 & w16412) | (~w7775 & w16412);
assign w7963 = (w7199 & ~w7727) | (w7199 & w16413) | (~w7727 & w16413);
assign w7964 = (w6999 & w17668) | (w6999 & ~w7647) | (w17668 & ~w7647);
assign w7965 = ~w6195 & ~w7860;
assign w7966 = w7180 & w7965;
assign w7967 = w7884 & w16414;
assign w7968 = (w7185 & ~w16414) | (w7185 & w17199) | (~w16414 & w17199);
assign w7969 = (w7188 & ~w7854) | (w7188 & w17669) | (~w7854 & w17669);
assign w7970 = (w7176 & ~w7695) | (w7176 & w17200) | (~w7695 & w17200);
assign w7971 = ~w7957 & ~w7961;
assign w7972 = ~w7962 & ~w7963;
assign w7973 = ~w7964 & ~w7968;
assign w7974 = ~w7969 & ~w7970;
assign w7975 = w7973 & w7974;
assign w7976 = w7971 & w7972;
assign w7977 = w7975 & w7976;
assign w7978 = (w7167 & ~w7826) | (w7167 & w17201) | (~w7826 & w17201);
assign w7979 = (w7214 & ~w7228) | (w7214 & w18062) | (~w7228 & w18062);
assign w7980 = (w7164 & ~w7601) | (w7164 & w16415) | (~w7601 & w16415);
assign w7981 = (w7168 & ~w7210) | (w7168 & w17202) | (~w7210 & w17202);
assign w7982 = w7087 & ~w7585;
assign w7983 = (w7193 & ~w7623) | (w7193 & w16416) | (~w7623 & w16416);
assign w7984 = w7058 & ~w7982;
assign w7985 = ~w7979 & w7984;
assign w7986 = ~w7980 & ~w7983;
assign w7987 = w7985 & w7986;
assign w7988 = ~w7978 & w7981;
assign w7989 = w7987 & w7988;
assign w7990 = w7977 & w7989;
assign w7991 = pi017 & w7990;
assign w7992 = w7646 & w18330;
assign w7993 = w7347 & ~w7585;
assign w7994 = ~w5679 & ~w6962;
assign w7995 = ~w7027 & w7994;
assign w7996 = ~w6935 & w7536;
assign w7997 = ~w4867 & ~w5652;
assign w7998 = ~w1980 & ~w3533;
assign w7999 = ~w4581 & w7998;
assign w8000 = w7997 & w7999;
assign w8001 = ~w2903 & ~w4725;
assign w8002 = w8000 & w8001;
assign w8003 = ~pi199 & pi207;
assign w8004 = pi199 & ~pi207;
assign w8005 = ~pi200 & pi208;
assign w8006 = pi200 & ~pi208;
assign w8007 = ~pi201 & pi209;
assign w8008 = pi201 & ~pi209;
assign w8009 = pi202 & ~pi210;
assign w8010 = ~pi203 & pi211;
assign w8011 = ~pi202 & pi210;
assign w8012 = pi203 & ~pi211;
assign w8013 = pi204 & ~pi212;
assign w8014 = ~pi204 & pi212;
assign w8015 = pi205 & ~pi213;
assign w8016 = ~pi205 & pi213;
assign w8017 = pi206 & ~pi214;
assign w8018 = ~w8016 & w8017;
assign w8019 = ~w8015 & ~w8018;
assign w8020 = ~w8014 & ~w8019;
assign w8021 = ~w8012 & ~w8013;
assign w8022 = ~w8020 & w8021;
assign w8023 = ~w8010 & ~w8011;
assign w8024 = ~w8022 & w8023;
assign w8025 = ~w8008 & ~w8009;
assign w8026 = ~w8024 & w8025;
assign w8027 = ~w8007 & ~w8026;
assign w8028 = ~w8006 & ~w8027;
assign w8029 = ~w8005 & ~w8028;
assign w8030 = ~w8004 & ~w8029;
assign w8031 = ~w8003 & ~w8030;
assign w8032 = w6105 & ~w7565;
assign w8033 = ~w4894 & ~w6097;
assign w8034 = w8031 & w8033;
assign w8035 = w8032 & w8034;
assign w8036 = ~w2930 & ~w3532;
assign w8037 = ~w4608 & w8036;
assign w8038 = w1979 & w8037;
assign w8039 = ~w823 & w8002;
assign w8040 = ~w217 & w8039;
assign w8041 = w4729 & w8040;
assign w8042 = w7996 & w8041;
assign w8043 = w1755 & w8042;
assign w8044 = w6102 & w8043;
assign w8045 = w6101 & w8038;
assign w8046 = w8044 & w8045;
assign w8047 = w7995 & w8046;
assign w8048 = w8035 & w8047;
assign w8049 = ~w7000 & w8048;
assign w8050 = ~w7993 & w8049;
assign w8051 = w7992 & w8050;
assign w8052 = pi022 & w8051;
assign w8053 = ~w174 & w178;
assign w8054 = ~w170 & w8053;
assign w8055 = w184 & ~w8054;
assign w8056 = ~pi199 & pi271;
assign w8057 = pi199 & ~pi271;
assign w8058 = ~pi200 & pi272;
assign w8059 = pi200 & ~pi272;
assign w8060 = ~pi201 & pi273;
assign w8061 = pi201 & ~pi273;
assign w8062 = pi202 & ~pi274;
assign w8063 = ~pi203 & pi275;
assign w8064 = ~pi202 & pi274;
assign w8065 = pi203 & ~pi275;
assign w8066 = pi204 & ~pi276;
assign w8067 = ~pi204 & pi276;
assign w8068 = pi205 & ~pi277;
assign w8069 = ~pi205 & pi277;
assign w8070 = pi206 & ~pi278;
assign w8071 = ~w8069 & w8070;
assign w8072 = ~w8068 & ~w8071;
assign w8073 = ~w8067 & ~w8072;
assign w8074 = ~w8065 & ~w8066;
assign w8075 = ~w8073 & w8074;
assign w8076 = ~w8063 & ~w8064;
assign w8077 = ~w8075 & w8076;
assign w8078 = ~w8061 & ~w8062;
assign w8079 = ~w8077 & w8078;
assign w8080 = ~w8060 & ~w8079;
assign w8081 = ~w8059 & ~w8080;
assign w8082 = ~w8058 & ~w8081;
assign w8083 = ~w8057 & ~w8082;
assign w8084 = ~w8056 & ~w8083;
assign w8085 = pi199 & ~pi263;
assign w8086 = ~pi199 & pi263;
assign w8087 = pi200 & ~pi264;
assign w8088 = ~pi200 & pi264;
assign w8089 = pi201 & ~pi265;
assign w8090 = ~pi202 & pi266;
assign w8091 = ~pi201 & pi265;
assign w8092 = pi202 & ~pi266;
assign w8093 = ~pi203 & pi267;
assign w8094 = pi203 & ~pi267;
assign w8095 = ~pi204 & pi268;
assign w8096 = pi204 & ~pi268;
assign w8097 = ~pi205 & pi269;
assign w8098 = pi205 & ~pi269;
assign w8099 = pi206 & ~pi270;
assign w8100 = ~w8098 & ~w8099;
assign w8101 = ~w8097 & ~w8100;
assign w8102 = ~w8096 & ~w8101;
assign w8103 = ~w8095 & ~w8102;
assign w8104 = ~w8094 & ~w8103;
assign w8105 = ~w8093 & ~w8104;
assign w8106 = ~w8092 & ~w8105;
assign w8107 = ~w8090 & ~w8091;
assign w8108 = ~w8106 & w8107;
assign w8109 = ~w8089 & ~w8108;
assign w8110 = ~w8088 & ~w8109;
assign w8111 = ~w8087 & ~w8110;
assign w8112 = ~w8086 & ~w8111;
assign w8113 = ~w8085 & ~w8112;
assign w8114 = ~w8084 & w8113;
assign w8115 = ~pi199 & pi255;
assign w8116 = pi199 & ~pi255;
assign w8117 = ~pi200 & pi256;
assign w8118 = pi200 & ~pi256;
assign w8119 = ~pi201 & pi257;
assign w8120 = pi201 & ~pi257;
assign w8121 = pi202 & ~pi258;
assign w8122 = ~pi203 & pi259;
assign w8123 = ~pi202 & pi258;
assign w8124 = pi203 & ~pi259;
assign w8125 = pi204 & ~pi260;
assign w8126 = ~pi204 & pi260;
assign w8127 = pi205 & ~pi261;
assign w8128 = ~pi205 & pi261;
assign w8129 = pi206 & ~pi262;
assign w8130 = ~w8128 & w8129;
assign w8131 = ~w8127 & ~w8130;
assign w8132 = ~w8126 & ~w8131;
assign w8133 = ~w8124 & ~w8125;
assign w8134 = ~w8132 & w8133;
assign w8135 = ~w8122 & ~w8123;
assign w8136 = ~w8134 & w8135;
assign w8137 = ~w8120 & ~w8121;
assign w8138 = ~w8136 & w8137;
assign w8139 = ~w8119 & ~w8138;
assign w8140 = ~w8118 & ~w8139;
assign w8141 = ~w8117 & ~w8140;
assign w8142 = ~w8116 & ~w8141;
assign w8143 = ~w8115 & ~w8142;
assign w8144 = ~pi199 & pi247;
assign w8145 = pi199 & ~pi247;
assign w8146 = ~pi200 & pi248;
assign w8147 = pi200 & ~pi248;
assign w8148 = ~pi201 & pi249;
assign w8149 = pi201 & ~pi249;
assign w8150 = pi202 & ~pi250;
assign w8151 = ~pi203 & pi251;
assign w8152 = ~pi202 & pi250;
assign w8153 = pi203 & ~pi251;
assign w8154 = pi204 & ~pi252;
assign w8155 = ~pi204 & pi252;
assign w8156 = pi205 & ~pi253;
assign w8157 = ~pi205 & pi253;
assign w8158 = pi206 & ~pi254;
assign w8159 = ~w8157 & w8158;
assign w8160 = ~w8156 & ~w8159;
assign w8161 = ~w8155 & ~w8160;
assign w8162 = ~w8153 & ~w8154;
assign w8163 = ~w8161 & w8162;
assign w8164 = ~w8151 & ~w8152;
assign w8165 = ~w8163 & w8164;
assign w8166 = ~w8149 & ~w8150;
assign w8167 = ~w8165 & w8166;
assign w8168 = ~w8148 & ~w8167;
assign w8169 = ~w8147 & ~w8168;
assign w8170 = ~w8146 & ~w8169;
assign w8171 = ~w8145 & ~w8170;
assign w8172 = ~w8144 & ~w8171;
assign w8173 = ~w8143 & ~w8172;
assign w8174 = w8114 & w8173;
assign w8175 = ~pi199 & pi215;
assign w8176 = pi199 & ~pi215;
assign w8177 = ~pi200 & pi216;
assign w8178 = pi200 & ~pi216;
assign w8179 = ~pi201 & pi217;
assign w8180 = pi202 & ~pi218;
assign w8181 = pi201 & ~pi217;
assign w8182 = ~pi202 & pi218;
assign w8183 = pi203 & ~pi219;
assign w8184 = ~pi203 & pi219;
assign w8185 = pi204 & ~pi220;
assign w8186 = ~pi204 & pi220;
assign w8187 = ~pi205 & pi221;
assign w8188 = pi206 & ~pi222;
assign w8189 = ~w8187 & w8188;
assign w8190 = pi205 & ~pi221;
assign w8191 = ~w8189 & ~w8190;
assign w8192 = ~w8186 & ~w8191;
assign w8193 = ~w8185 & ~w8192;
assign w8194 = ~w8184 & ~w8193;
assign w8195 = ~w8183 & ~w8194;
assign w8196 = ~w8182 & ~w8195;
assign w8197 = ~w8180 & ~w8181;
assign w8198 = ~w8196 & w8197;
assign w8199 = ~w8179 & ~w8198;
assign w8200 = ~w8178 & ~w8199;
assign w8201 = ~w8177 & ~w8200;
assign w8202 = ~w8176 & ~w8201;
assign w8203 = ~w8175 & ~w8202;
assign w8204 = ~pi199 & pi239;
assign w8205 = pi199 & ~pi239;
assign w8206 = ~pi200 & pi240;
assign w8207 = pi200 & ~pi240;
assign w8208 = ~pi201 & pi241;
assign w8209 = pi201 & ~pi241;
assign w8210 = pi202 & ~pi242;
assign w8211 = ~pi203 & pi243;
assign w8212 = ~pi202 & pi242;
assign w8213 = pi203 & ~pi243;
assign w8214 = pi204 & ~pi244;
assign w8215 = ~pi204 & pi244;
assign w8216 = pi205 & ~pi245;
assign w8217 = ~pi205 & pi245;
assign w8218 = pi206 & ~pi246;
assign w8219 = ~w8217 & w8218;
assign w8220 = ~w8216 & ~w8219;
assign w8221 = ~w8215 & ~w8220;
assign w8222 = ~w8213 & ~w8214;
assign w8223 = ~w8221 & w8222;
assign w8224 = ~w8211 & ~w8212;
assign w8225 = ~w8223 & w8224;
assign w8226 = ~w8209 & ~w8210;
assign w8227 = ~w8225 & w8226;
assign w8228 = ~w8208 & ~w8227;
assign w8229 = ~w8207 & ~w8228;
assign w8230 = ~w8206 & ~w8229;
assign w8231 = ~w8205 & ~w8230;
assign w8232 = ~w8204 & ~w8231;
assign w8233 = pi199 & ~pi231;
assign w8234 = ~pi199 & pi231;
assign w8235 = pi200 & ~pi232;
assign w8236 = ~pi200 & pi232;
assign w8237 = pi201 & ~pi233;
assign w8238 = ~pi202 & pi234;
assign w8239 = ~pi201 & pi233;
assign w8240 = pi202 & ~pi234;
assign w8241 = ~pi203 & pi235;
assign w8242 = pi203 & ~pi235;
assign w8243 = ~pi204 & pi236;
assign w8244 = pi204 & ~pi236;
assign w8245 = ~pi205 & pi237;
assign w8246 = pi205 & ~pi237;
assign w8247 = pi206 & ~pi238;
assign w8248 = ~w8246 & ~w8247;
assign w8249 = ~w8245 & ~w8248;
assign w8250 = ~w8244 & ~w8249;
assign w8251 = ~w8243 & ~w8250;
assign w8252 = ~w8242 & ~w8251;
assign w8253 = ~w8241 & ~w8252;
assign w8254 = ~w8240 & ~w8253;
assign w8255 = ~w8238 & ~w8239;
assign w8256 = ~w8254 & w8255;
assign w8257 = ~w8237 & ~w8256;
assign w8258 = ~w8236 & ~w8257;
assign w8259 = ~w8235 & ~w8258;
assign w8260 = ~w8234 & ~w8259;
assign w8261 = ~w8233 & ~w8260;
assign w8262 = ~w8232 & w8261;
assign w8263 = pi199 & ~pi223;
assign w8264 = ~pi199 & pi223;
assign w8265 = pi200 & ~pi224;
assign w8266 = ~pi200 & pi224;
assign w8267 = pi201 & ~pi225;
assign w8268 = ~pi201 & pi225;
assign w8269 = pi202 & ~pi226;
assign w8270 = ~pi202 & pi226;
assign w8271 = pi203 & ~pi227;
assign w8272 = ~pi203 & pi227;
assign w8273 = ~pi204 & pi228;
assign w8274 = pi205 & ~pi229;
assign w8275 = ~pi205 & pi229;
assign w8276 = pi206 & ~pi230;
assign w8277 = ~w8275 & w8276;
assign w8278 = ~w8274 & ~w8277;
assign w8279 = ~w8273 & ~w8278;
assign w8280 = pi204 & ~pi228;
assign w8281 = ~w8279 & ~w8280;
assign w8282 = ~w8272 & ~w8281;
assign w8283 = ~w8271 & ~w8282;
assign w8284 = ~w8270 & ~w8283;
assign w8285 = ~w8269 & ~w8284;
assign w8286 = ~w8268 & ~w8285;
assign w8287 = ~w8267 & ~w8286;
assign w8288 = ~w8266 & ~w8287;
assign w8289 = ~w8265 & ~w8288;
assign w8290 = ~w8264 & ~w8289;
assign w8291 = ~w8263 & ~w8290;
assign w8292 = ~w8203 & w8262;
assign w8293 = w8291 & w8292;
assign w8294 = w8174 & w8293;
assign w8295 = pi135 & w4714;
assign w8296 = w7529 & w8295;
assign w8297 = pi039 & w8296;
assign w8298 = ~pi199 & w4726;
assign w8299 = ~w8297 & ~w8298;
assign w8300 = w2627 & w4717;
assign w8301 = w6965 & w8300;
assign w8302 = ~w2009 & ~w8299;
assign w8303 = ~w8055 & w8302;
assign w8304 = ~w1727 & w8303;
assign w8305 = ~w2901 & ~w3504;
assign w8306 = ~w4637 & ~w5737;
assign w8307 = ~w7056 & w7996;
assign w8308 = w8306 & w8307;
assign w8309 = w8304 & w8305;
assign w8310 = w4062 & w7566;
assign w8311 = w8309 & w8310;
assign w8312 = w8308 & w8311;
assign w8313 = ~w7259 & w8301;
assign w8314 = w8312 & w8313;
assign w8315 = ~w8031 & w8314;
assign w8316 = w8032 & w8315;
assign w8317 = w8294 & w8316;
assign w8318 = ~w4923 & w8317;
assign w8319 = w7992 & w8318;
assign w8320 = pi021 & w8319;
assign w8321 = (w7215 & ~w16414) | (w7215 & w17203) | (~w16414 & w17203);
assign w8322 = (w7219 & ~w7775) | (w7219 & w16417) | (~w7775 & w16417);
assign w8323 = ~w8321 & ~w8322;
assign w8324 = (w7220 & ~w7826) | (w7220 & w17204) | (~w7826 & w17204);
assign w8325 = (w7213 & ~w7727) | (w7213 & w16418) | (~w7727 & w16418);
assign w8326 = w7186 & ~w7750;
assign w8327 = (w7225 & ~w7695) | (w7225 & w17205) | (~w7695 & w17205);
assign w8328 = (w7223 & ~w7854) | (w7223 & w17670) | (~w7854 & w17670);
assign w8329 = (w7224 & ~w7919) | (w7224 & w17671) | (~w7919 & w17671);
assign w8330 = w7979 & ~w8326;
assign w8331 = ~w8327 & w8330;
assign w8332 = ~w8328 & ~w8329;
assign w8333 = w8331 & w8332;
assign w8334 = ~w8324 & ~w8325;
assign w8335 = w8323 & w8334;
assign w8336 = w8333 & w8335;
assign w8337 = pi014 & w8336;
assign w8338 = w7594 & ~w7960;
assign w8339 = (w7587 & ~w7775) | (w7587 & w16419) | (~w7775 & w16419);
assign w8340 = (w7166 & ~w7826) | (w7166 & w17206) | (~w7826 & w17206);
assign w8341 = ~w2695 & w8340;
assign w8342 = (w7222 & ~w7854) | (w7222 & w17672) | (~w7854 & w17672);
assign w8343 = ~w2444 & w8342;
assign w8344 = (w7175 & ~w7695) | (w7175 & w17207) | (~w7695 & w17207);
assign w8345 = ~w5224 & w8344;
assign w8346 = w7593 & ~w7701;
assign w8347 = w7184 & ~w7967;
assign w8348 = w691 & w8347;
assign w8349 = (w7588 & ~w7727) | (w7588 & w18331) | (~w7727 & w18331);
assign w8350 = ~w7979 & w7980;
assign w8351 = ~w8338 & w8350;
assign w8352 = ~w8339 & ~w8346;
assign w8353 = ~w8349 & w8352;
assign w8354 = ~w8341 & w8351;
assign w8355 = ~w8343 & ~w8345;
assign w8356 = ~w8348 & w8355;
assign w8357 = w8353 & w8354;
assign w8358 = w8356 & w8357;
assign w8359 = pi016 & w8358;
assign w8360 = (w7632 & ~w7695) | (w7632 & w17208) | (~w7695 & w17208);
assign w8361 = (w7636 & ~w7775) | (w7636 & w16420) | (~w7775 & w16420);
assign w8362 = (~w6447 & ~w7663) | (~w6447 & w17673) | (~w7663 & w17673);
assign w8363 = w7633 & w8362;
assign w8364 = (w7638 & ~w7826) | (w7638 & w17209) | (~w7826 & w17209);
assign w8365 = (w7639 & ~w7854) | (w7639 & w17674) | (~w7854 & w17674);
assign w8366 = w7626 & ~w7967;
assign w8367 = (w7630 & ~w7210) | (w7630 & w18063) | (~w7210 & w18063);
assign w8368 = (~w7192 & ~w7623) | (~w7192 & w16421) | (~w7623 & w16421);
assign w8369 = w7565 & ~w7585;
assign w8370 = w7637 & ~w7960;
assign w8371 = (w7629 & ~w7727) | (w7629 & w17675) | (~w7727 & w17675);
assign w8372 = (~w8369 & w17676) | (~w8369 & ~w7647) | (w17676 & ~w7647);
assign w8373 = ~w8368 & w8372;
assign w8374 = ~w8360 & ~w8361;
assign w8375 = ~w8364 & ~w8365;
assign w8376 = ~w8366 & ~w8367;
assign w8377 = ~w8370 & ~w8371;
assign w8378 = w8376 & w8377;
assign w8379 = w8374 & w8375;
assign w8380 = ~w8363 & w8373;
assign w8381 = w8379 & w8380;
assign w8382 = w8378 & w8381;
assign w8383 = pi020 & w8382;
assign w8384 = (w7611 & ~w7695) | (w7611 & w17210) | (~w7695 & w17210);
assign w8385 = w2416 & w8342;
assign w8386 = ~w7980 & w8368;
assign w8387 = ~w8384 & w8386;
assign w8388 = ~w8385 & w8387;
assign w8389 = (w7196 & ~w7775) | (w7196 & w16422) | (~w7775 & w16422);
assign w8390 = ~w3623 & w8389;
assign w8391 = w7607 & ~w7701;
assign w8392 = (w7606 & ~w7210) | (w7606 & w18064) | (~w7210 & w18064);
assign w8393 = (w7608 & ~w7826) | (w7608 & w18065) | (~w7826 & w18065);
assign w8394 = (w7613 & ~w16414) | (w7613 & w17211) | (~w16414 & w17211);
assign w8395 = (w7609 & ~w7919) | (w7609 & w17677) | (~w7919 & w17677);
assign w8396 = (w7610 & ~w7727) | (w7610 & w17678) | (~w7727 & w17678);
assign w8397 = ~w8392 & ~w8393;
assign w8398 = ~w8394 & ~w8395;
assign w8399 = ~w8396 & w8398;
assign w8400 = w8397 & w8399;
assign w8401 = ~w8390 & ~w8391;
assign w8402 = w8388 & w8401;
assign w8403 = w8400 & w8402;
assign w8404 = pi018 & w8403;
assign w8405 = ~w3949 & w8389;
assign w8406 = (~w7565 & w17679) | (~w7565 & ~w7647) | (w17679 & ~w7647);
assign w8407 = w7528 & ~w7585;
assign w8408 = ~w6128 & w7656;
assign w8409 = (w8408 & ~w7663) | (w8408 & w17680) | (~w7663 & w17680);
assign w8410 = ~w821 & w7184;
assign w8411 = (w8410 & ~w16414) | (w8410 & w17212) | (~w16414 & w17212);
assign w8412 = w1668 & w7173;
assign w8413 = (w8412 & ~w7919) | (w8412 & w17681) | (~w7919 & w17681);
assign w8414 = ~w4551 & w7198;
assign w8415 = (w8414 & ~w7727) | (w8414 & w16423) | (~w7727 & w16423);
assign w8416 = (w17206 & w17682) | (w17206 & w17683) | (w17682 & w17683);
assign w8417 = (~w7695 & w18066) | (~w7695 & w18067) | (w18066 & w18067);
assign w8418 = (~w7113 & ~w7210) | (~w7113 & w17213) | (~w7210 & w17213);
assign w8419 = (~w7210 & w18068) | (~w7210 & w18069) | (w18068 & w18069);
assign w8420 = ~w2042 & w8342;
assign w8421 = w7349 & w8407;
assign w8422 = ~w8368 & w8421;
assign w8423 = ~w8406 & w8422;
assign w8424 = ~w8409 & ~w8411;
assign w8425 = ~w8413 & ~w8415;
assign w8426 = w8424 & w8425;
assign w8427 = ~w8405 & w8423;
assign w8428 = ~w8416 & ~w8417;
assign w8429 = ~w8419 & ~w8420;
assign w8430 = w8428 & w8429;
assign w8431 = w8426 & w8427;
assign w8432 = w8430 & w8431;
assign w8433 = pi019 & w8432;
assign w8434 = (w7654 & ~w7826) | (w7654 & w17214) | (~w7826 & w17214);
assign w8435 = w5828 & ~w7585;
assign w8436 = w5740 & ~w6447;
assign w8437 = ~w8435 & w8436;
assign w8438 = (w8437 & ~w7663) | (w8437 & w17684) | (~w7663 & w17684);
assign w8439 = ~w8434 & w8438;
assign w8440 = (w16415 & w17215) | (w16415 & w17216) | (w17215 & w17216);
assign w8441 = (w7651 & ~w7695) | (w7651 & w17217) | (~w7695 & w17217);
assign w8442 = (w7665 & ~w7854) | (w7665 & w17685) | (~w7854 & w17685);
assign w8443 = (~w5769 & w17686) | (~w5769 & ~w7647) | (w17686 & ~w7647);
assign w8444 = (w7652 & ~w16414) | (w7652 & w17218) | (~w16414 & w17218);
assign w8445 = (w7667 & ~w7775) | (w7667 & w17687) | (~w7775 & w17687);
assign w8446 = ~w7979 & ~w8440;
assign w8447 = ~w8441 & ~w8442;
assign w8448 = ~w8443 & ~w8444;
assign w8449 = ~w8445 & w8448;
assign w8450 = w8446 & w8447;
assign w8451 = w8449 & w8450;
assign w8452 = (w7664 & ~w7919) | (w7664 & w17688) | (~w7919 & w17688);
assign w8453 = w5857 & w8368;
assign w8454 = (w7655 & ~w7210) | (w7655 & w17219) | (~w7210 & w17219);
assign w8455 = (w7650 & ~w7727) | (w7650 & w16424) | (~w7727 & w16424);
assign w8456 = ~w8452 & ~w8453;
assign w8457 = ~w8454 & ~w8455;
assign w8458 = w8456 & w8457;
assign w8459 = w8451 & w8458;
assign w8460 = w8439 & w8459;
assign w8461 = w6376 & w8460;
assign w8462 = w4984 & w8344;
assign w8463 = w5163 & w8462;
assign w8464 = ~pi013 & w8463;
assign w8465 = ~w5192 & ~w7585;
assign w8466 = (w7677 & ~w7775) | (w7677 & w18332) | (~w7775 & w18332);
assign w8467 = w4925 & ~w8465;
assign w8468 = ~w8466 & w8467;
assign w8469 = ~w8326 & w8468;
assign w8470 = w7173 & ~w7960;
assign w8471 = ~w7960 & w18333;
assign w8472 = (w7683 & ~w7601) | (w7683 & w16425) | (~w7601 & w16425);
assign w8473 = (w7674 & ~w7228) | (w7674 & w18070) | (~w7228 & w18070);
assign w8474 = w5341 & w8368;
assign w8475 = w5282 & ~w7648;
assign w8476 = (w7676 & ~w7826) | (w7676 & w17220) | (~w7826 & w17220);
assign w8477 = w7681 & ~w7967;
assign w8478 = w7680 & ~w7701;
assign w8479 = (~w6523 & ~w7727) | (~w6523 & w16426) | (~w7727 & w16426);
assign w8480 = w6428 & w8479;
assign w8481 = (w7682 & ~w7854) | (w7682 & w18334) | (~w7854 & w18334);
assign w8482 = (w7678 & ~w7210) | (w7678 & w18335) | (~w7210 & w18335);
assign w8483 = ~w8472 & ~w8473;
assign w8484 = ~w8474 & w8483;
assign w8485 = ~w8475 & ~w8476;
assign w8486 = ~w8477 & ~w8478;
assign w8487 = ~w8481 & ~w8482;
assign w8488 = w8486 & w8487;
assign w8489 = w8484 & w8485;
assign w8490 = ~w8471 & ~w8480;
assign w8491 = w8489 & w8490;
assign w8492 = w8488 & w8491;
assign w8493 = w8469 & w8492;
assign w8494 = w8464 & w8493;
assign w8495 = ~w8434 & w17689;
assign w8496 = w8458 & w8495;
assign w8497 = w8451 & w8496;
assign w8498 = ~w8336 & ~w8497;
assign w8499 = (w7705 & ~w17182) | (w7705 & w17690) | (~w17182 & w17690);
assign w8500 = (w7743 & ~w7919) | (w7743 & w17691) | (~w7919 & w17691);
assign w8501 = (w7742 & ~w7775) | (w7742 & w16427) | (~w7775 & w16427);
assign w8502 = (w7741 & ~w16414) | (w7741 & w17221) | (~w16414 & w17221);
assign w8503 = (w7737 & ~w7727) | (w7737 & w16428) | (~w7727 & w16428);
assign w8504 = (w7738 & ~w7826) | (w7738 & w17222) | (~w7826 & w17222);
assign w8505 = (w7740 & ~w7854) | (w7740 & w18336) | (~w7854 & w18336);
assign w8506 = w8326 & ~w8499;
assign w8507 = ~w8500 & w8506;
assign w8508 = ~w8501 & ~w8502;
assign w8509 = ~w8503 & ~w8504;
assign w8510 = ~w8505 & w8509;
assign w8511 = w8507 & w8508;
assign w8512 = w8510 & w8511;
assign w8513 = pi012 & w8512;
assign w8514 = ~w5431 & w8463;
assign w8515 = w8469 & w8514;
assign w8516 = w8492 & w8515;
assign w8517 = ~w7603 & w7713;
assign w8518 = w7706 & ~w7960;
assign w8519 = (w7703 & ~w7210) | (w7703 & w18071) | (~w7210 & w18071);
assign w8520 = ~w7701 & w7719;
assign w8521 = w7715 & ~w7967;
assign w8522 = (w7716 & ~w7775) | (w7716 & w16429) | (~w7775 & w16429);
assign w8523 = (w7717 & ~w7826) | (w7717 & w18072) | (~w7826 & w18072);
assign w8524 = (w7714 & ~w7854) | (w7714 & w18073) | (~w7854 & w18073);
assign w8525 = (w7704 & ~w7750) | (w7704 & w18337) | (~w7750 & w18337);
assign w8526 = (w7720 & ~w7695) | (w7720 & w18074) | (~w7695 & w18074);
assign w8527 = ~w4371 & ~w7648;
assign w8528 = w4163 & w7979;
assign w8529 = w4551 & ~w7585;
assign w8530 = ~w4400 & w8368;
assign w8531 = ~w8499 & ~w8529;
assign w8532 = ~w8517 & w8531;
assign w8533 = w8479 & ~w8518;
assign w8534 = ~w8519 & ~w8520;
assign w8535 = ~w8521 & ~w8522;
assign w8536 = ~w8523 & ~w8524;
assign w8537 = ~w8525 & ~w8526;
assign w8538 = ~w8527 & ~w8528;
assign w8539 = ~w8530 & w8538;
assign w8540 = w8536 & w8537;
assign w8541 = w8534 & w8535;
assign w8542 = w8532 & w8533;
assign w8543 = w8541 & w8542;
assign w8544 = w8539 & w8540;
assign w8545 = w8543 & w8544;
assign w8546 = w7712 & w8545;
assign w8547 = w7735 & w8546;
assign w8548 = w6521 & w8545;
assign w8549 = ~w3254 & ~w3296;
assign w8550 = ~w4705 & w8549;
assign w8551 = ~w6219 & w8550;
assign w8552 = ~pi007 & w8551;
assign w8553 = (w7800 & ~w7775) | (w7800 & w16430) | (~w7775 & w16430);
assign w8554 = (w7801 & ~w7663) | (w7801 & w17692) | (~w7663 & w17692);
assign w8555 = ~w8553 & ~w8554;
assign w8556 = w2932 & w3019;
assign w8557 = (~w8556 & ~w7647) | (~w8556 & w17693) | (~w7647 & w17693);
assign w8558 = w3225 & ~w7585;
assign w8559 = ~w7750 & w7814;
assign w8560 = (w7809 & ~w7854) | (w7809 & w17694) | (~w7854 & w17694);
assign w8561 = (w7812 & ~w7727) | (w7812 & w16431) | (~w7727 & w16431);
assign w8562 = ~w5431 & w7798;
assign w8563 = ~w6558 & w8562;
assign w8564 = (w8563 & ~w7826) | (w8563 & w17223) | (~w7826 & w17223);
assign w8565 = (~w8558 & w7750) | (~w8558 & w17695) | (w7750 & w17695);
assign w8566 = ~w8560 & w8565;
assign w8567 = ~w8561 & w8564;
assign w8568 = w8566 & w8567;
assign w8569 = (w7805 & ~w16414) | (w7805 & w17224) | (~w16414 & w17224);
assign w8570 = (w7810 & ~w7228) | (w7810 & w18075) | (~w7228 & w18075);
assign w8571 = (w7799 & ~w7919) | (w7799 & w17696) | (~w7919 & w17696);
assign w8572 = (w7813 & ~w7210) | (w7813 & w17225) | (~w7210 & w17225);
assign w8573 = (w16415 & w17226) | (w16415 & w17227) | (w17226 & w17227);
assign w8574 = (w7808 & ~w7695) | (w7808 & w17228) | (~w7695 & w17228);
assign w8575 = w2723 & w8368;
assign w8576 = ~w8569 & ~w8570;
assign w8577 = ~w8571 & ~w8572;
assign w8578 = ~w8573 & ~w8574;
assign w8579 = ~w8575 & w8578;
assign w8580 = w8576 & w8577;
assign w8581 = w8579 & w8580;
assign w8582 = w8555 & ~w8557;
assign w8583 = w8568 & w8582;
assign w8584 = w8581 & w8583;
assign w8585 = ~w3402 & w5524;
assign w8586 = ~w5531 & w8585;
assign w8587 = w8584 & w8586;
assign w8588 = w8552 & w8587;
assign w8589 = (w7761 & ~w7826) | (w7761 & w18338) | (~w7826 & w18338);
assign w8590 = ~w3773 & w3919;
assign w8591 = w7196 & w8590;
assign w8592 = (w8591 & ~w7775) | (w8591 & w16432) | (~w7775 & w16432);
assign w8593 = w3831 & w8592;
assign w8594 = (w7762 & ~w7601) | (w7762 & w16433) | (~w7601 & w16433);
assign w8595 = w3949 & ~w7584;
assign w8596 = (w7760 & ~w7663) | (w7760 & w17697) | (~w7663 & w17697);
assign w8597 = (w7756 & ~w7695) | (w7756 & w17229) | (~w7695 & w17229);
assign w8598 = (~w3565 & w17698) | (~w3565 & ~w7647) | (w17698 & ~w7647);
assign w8599 = w3536 & ~w8595;
assign w8600 = (~w16433 & w17230) | (~w16433 & w17231) | (w17230 & w17231);
assign w8601 = ~w8596 & w8600;
assign w8602 = ~w8597 & ~w8598;
assign w8603 = w8601 & w8602;
assign w8604 = (w7777 & ~w7727) | (w7777 & w16434) | (~w7727 & w16434);
assign w8605 = (w7755 & ~w7919) | (w7755 & w17699) | (~w7919 & w17699);
assign w8606 = (w7776 & ~w16414) | (w7776 & w17232) | (~w16414 & w17232);
assign w8607 = (~w7759 & ~w7750) | (~w7759 & w17700) | (~w7750 & w17700);
assign w8608 = (w7763 & ~w7854) | (w7763 & w17701) | (~w7854 & w17701);
assign w8609 = (w7764 & ~w7228) | (w7764 & w17884) | (~w7228 & w17884);
assign w8610 = (w7765 & ~w7623) | (w7765 & w16435) | (~w7623 & w16435);
assign w8611 = (w7766 & ~w7210) | (w7766 & w17885) | (~w7210 & w17885);
assign w8612 = ~w8609 & ~w8610;
assign w8613 = ~w8604 & w8612;
assign w8614 = ~w8605 & ~w8606;
assign w8615 = ~w8607 & ~w8608;
assign w8616 = ~w8611 & w8615;
assign w8617 = w8613 & w8614;
assign w8618 = w8616 & w8617;
assign w8619 = ~w8589 & w8593;
assign w8620 = w8603 & w8619;
assign w8621 = w8618 & w8620;
assign w8622 = (w7902 & ~w7775) | (w7902 & w16436) | (~w7775 & w16436);
assign w8623 = ~w1668 & ~w7585;
assign w8624 = (w7908 & ~w7623) | (w7908 & w16437) | (~w7623 & w16437);
assign w8625 = (w7904 & ~w7228) | (w7904 & w17886) | (~w7228 & w17886);
assign w8626 = (w7910 & ~w7601) | (w7910 & w16438) | (~w7601 & w16438);
assign w8627 = ~w7750 & w7923;
assign w8628 = (w7907 & ~w7854) | (w7907 & w17887) | (~w7854 & w17887);
assign w8629 = (w7905 & ~w7826) | (w7905 & w17888) | (~w7826 & w17888);
assign w8630 = (w1168 & w17889) | (w1168 & ~w7647) | (w17889 & ~w7647);
assign w8631 = (w7903 & ~w16414) | (w7903 & w17890) | (~w16414 & w17890);
assign w8632 = w6631 & w8362;
assign w8633 = (w7924 & ~w7727) | (w7924 & w16439) | (~w7727 & w16439);
assign w8634 = (w7922 & ~w7695) | (w7922 & w17891) | (~w7695 & w17891);
assign w8635 = (w7906 & ~w7210) | (w7906 & w18339) | (~w7210 & w18339);
assign w8636 = w1548 & w1641;
assign w8637 = ~w3346 & w8636;
assign w8638 = w6382 & w18477;
assign w8639 = w7921 & w8638;
assign w8640 = ~w8623 & w8639;
assign w8641 = (w8640 & ~w7919) | (w8640 & w17892) | (~w7919 & w17892);
assign w8642 = ~w8624 & ~w8625;
assign w8643 = ~w8626 & ~w8627;
assign w8644 = w8642 & w8643;
assign w8645 = ~w8622 & w8641;
assign w8646 = ~w8628 & ~w8629;
assign w8647 = ~w8630 & ~w8631;
assign w8648 = ~w8633 & ~w8634;
assign w8649 = ~w8635 & w8648;
assign w8650 = w8646 & w8647;
assign w8651 = w8644 & w17893;
assign w8652 = w8649 & w8650;
assign w8653 = w8651 & w8652;
assign w8654 = w5565 & w8653;
assign w8655 = (w7647 & w18076) | (w7647 & w18077) | (w18076 & w18077);
assign w8656 = w8555 & w8655;
assign w8657 = w8568 & w8656;
assign w8658 = w8581 & w8657;
assign w8659 = (~w249 & w17702) | (~w249 & ~w7647) | (w17702 & ~w7647);
assign w8660 = (w821 & ~w7584) | (w821 & w17894) | (~w7584 & w17894);
assign w8661 = ~w7872 & w17895;
assign w8662 = ~w7750 & w7862;
assign w8663 = ~w8660 & w8661;
assign w8664 = (w8663 & ~w16414) | (w8663 & w17233) | (~w16414 & w17233);
assign w8665 = ~w8662 & w8664;
assign w8666 = (w7868 & ~w7695) | (w7868 & w17234) | (~w7695 & w17234);
assign w8667 = (w7870 & ~w7727) | (w7870 & w16440) | (~w7727 & w16440);
assign w8668 = (w7867 & ~w7854) | (w7867 & w17703) | (~w7854 & w17703);
assign w8669 = (w7871 & ~w7775) | (w7871 & w16441) | (~w7775 & w16441);
assign w8670 = (w7864 & ~w7919) | (w7864 & w17704) | (~w7919 & w17704);
assign w8671 = (w7860 & ~w7210) | (w7860 & w17896) | (~w7210 & w17896);
assign w8672 = (w7863 & ~w7228) | (w7863 & w17897) | (~w7228 & w17897);
assign w8673 = ~w8666 & ~w8672;
assign w8674 = ~w8667 & ~w8668;
assign w8675 = ~w8669 & ~w8670;
assign w8676 = ~w8671 & w8675;
assign w8677 = w8673 & w8674;
assign w8678 = w8676 & w8677;
assign w8679 = (w7869 & ~w7826) | (w7869 & w17235) | (~w7826 & w17235);
assign w8680 = (w7866 & ~w7601) | (w7866 & w16442) | (~w7601 & w16442);
assign w8681 = (w7865 & ~w7623) | (w7865 & w16443) | (~w7623 & w16443);
assign w8682 = (w7861 & ~w7663) | (w7861 & w17705) | (~w7663 & w17705);
assign w8683 = ~w8680 & ~w8681;
assign w8684 = w8683 & w17236;
assign w8685 = ~w7183 & ~w8659;
assign w8686 = w8665 & w8685;
assign w8687 = w8684 & w8686;
assign w8688 = w8678 & w8687;
assign w8689 = w7894 & w8688;
assign w8690 = (w7847 & ~w16414) | (w7847 & w17237) | (~w16414 & w17237);
assign w8691 = (w7840 & ~w7919) | (w7840 & w17706) | (~w7919 & w17706);
assign w8692 = (w7829 & ~w7210) | (w7829 & w17238) | (~w7210 & w17238);
assign w8693 = (w7846 & ~w7727) | (w7846 & w16444) | (~w7727 & w16444);
assign w8694 = (w16415 & w17239) | (w16415 & w17240) | (w17239 & w17240);
assign w8695 = (w7835 & ~w7623) | (w7835 & w16445) | (~w7623 & w16445);
assign w8696 = w2042 & ~w7585;
assign w8697 = w7221 & w7226;
assign w8698 = (w7844 & ~w7218) | (w7844 & w17707) | (~w7218 & w17707);
assign w8699 = ~w7750 & w7834;
assign w8700 = (w7841 & ~w7695) | (w7841 & w17241) | (~w7695 & w17241);
assign w8701 = w2012 & w7832;
assign w8702 = ~w8696 & w8701;
assign w8703 = ~w8695 & w8702;
assign w8704 = ~w8698 & ~w8699;
assign w8705 = w8703 & w8704;
assign w8706 = ~w8690 & ~w8691;
assign w8707 = ~w8692 & ~w8693;
assign w8708 = ~w8694 & ~w8700;
assign w8709 = w8707 & w8708;
assign w8710 = w8705 & w8706;
assign w8711 = w8709 & w8710;
assign w8712 = (w7843 & ~w7826) | (w7843 & w17898) | (~w7826 & w17898);
assign w8713 = (w7839 & ~w7854) | (w7839 & w17708) | (~w7854 & w17708);
assign w8714 = w6621 & w6663;
assign w8715 = w8714 & w8713;
assign w8716 = (~w2322 & w17709) | (~w2322 & ~w7647) | (w17709 & ~w7647);
assign w8717 = (w7845 & ~w7775) | (w7845 & w16446) | (~w7775 & w16446);
assign w8718 = (w7833 & ~w7663) | (w7833 & w17899) | (~w7663 & w17899);
assign w8719 = ~w8716 & ~w8717;
assign w8720 = ~w8718 & w8719;
assign w8721 = ~w8712 & w8715;
assign w8722 = w8720 & w8721;
assign w8723 = w8711 & w8722;
assign w8724 = pi005 & w8723;
assign w8725 = ~w8654 & ~w8658;
assign w8726 = ~w8689 & ~w8724;
assign w8727 = w8725 & w8726;
assign w8728 = ~w8588 & ~w8621;
assign w8729 = ~w8727 & w8728;
assign w8730 = pi009 & w8621;
assign w8731 = ~w8548 & ~w8730;
assign w8732 = ~w8729 & w8731;
assign w8733 = ~w8512 & ~w8547;
assign w8734 = ~w8732 & w8733;
assign w8735 = ~w8513 & ~w8516;
assign w8736 = ~w8734 & w8735;
assign w8737 = ~w8494 & w8498;
assign w8738 = ~w8736 & w8737;
assign w8739 = ~w8052 & ~w8320;
assign w8740 = ~w8337 & w8739;
assign w8741 = ~w7991 & w8740;
assign w8742 = ~w8359 & ~w8383;
assign w8743 = ~w8404 & ~w8433;
assign w8744 = w8742 & w8743;
assign w8745 = ~w8461 & w8741;
assign w8746 = w8744 & w8745;
assign w8747 = ~w8738 & w8746;
assign w8748 = ~w1729 & w2549;
assign w8749 = pi216 & ~pi256;
assign w8750 = ~pi216 & pi256;
assign w8751 = pi217 & ~pi257;
assign w8752 = ~pi217 & pi257;
assign w8753 = pi218 & ~pi258;
assign w8754 = ~pi219 & pi259;
assign w8755 = ~pi218 & pi258;
assign w8756 = pi219 & ~pi259;
assign w8757 = pi220 & ~pi260;
assign w8758 = ~pi220 & pi260;
assign w8759 = pi221 & ~pi261;
assign w8760 = ~pi221 & pi261;
assign w8761 = pi222 & ~pi262;
assign w8762 = ~w8760 & w8761;
assign w8763 = ~w8759 & ~w8762;
assign w8764 = ~w8758 & ~w8763;
assign w8765 = ~w8756 & ~w8757;
assign w8766 = ~w8764 & w8765;
assign w8767 = ~w8754 & ~w8755;
assign w8768 = ~w8766 & w8767;
assign w8769 = ~w8753 & ~w8768;
assign w8770 = ~w8752 & ~w8769;
assign w8771 = ~w8751 & ~w8770;
assign w8772 = ~w8750 & ~w8771;
assign w8773 = ~w8749 & ~w8772;
assign w8774 = pi215 & ~w8773;
assign w8775 = pi255 & ~w8774;
assign w8776 = ~pi215 & w8773;
assign w8777 = ~w8775 & ~w8776;
assign w8778 = ~pi215 & pi271;
assign w8779 = pi215 & ~pi271;
assign w8780 = ~pi216 & pi272;
assign w8781 = pi216 & ~pi272;
assign w8782 = ~pi217 & pi273;
assign w8783 = pi217 & ~pi273;
assign w8784 = pi218 & ~pi274;
assign w8785 = ~pi219 & pi275;
assign w8786 = ~pi218 & pi274;
assign w8787 = pi219 & ~pi275;
assign w8788 = pi220 & ~pi276;
assign w8789 = ~pi220 & pi276;
assign w8790 = pi221 & ~pi277;
assign w8791 = ~pi221 & pi277;
assign w8792 = pi222 & ~pi278;
assign w8793 = ~w8791 & w8792;
assign w8794 = ~w8790 & ~w8793;
assign w8795 = ~w8789 & ~w8794;
assign w8796 = ~w8787 & ~w8788;
assign w8797 = ~w8795 & w8796;
assign w8798 = ~w8785 & ~w8786;
assign w8799 = ~w8797 & w8798;
assign w8800 = ~w8783 & ~w8784;
assign w8801 = ~w8799 & w8800;
assign w8802 = ~w8782 & ~w8801;
assign w8803 = ~w8781 & ~w8802;
assign w8804 = ~w8780 & ~w8803;
assign w8805 = ~w8779 & ~w8804;
assign w8806 = ~w8778 & ~w8805;
assign w8807 = ~pi215 & pi263;
assign w8808 = pi215 & ~pi263;
assign w8809 = ~pi216 & pi264;
assign w8810 = pi216 & ~pi264;
assign w8811 = ~pi217 & pi265;
assign w8812 = pi217 & ~pi265;
assign w8813 = pi218 & ~pi266;
assign w8814 = ~pi219 & pi267;
assign w8815 = ~pi218 & pi266;
assign w8816 = pi219 & ~pi267;
assign w8817 = pi220 & ~pi268;
assign w8818 = ~pi220 & pi268;
assign w8819 = pi221 & ~pi269;
assign w8820 = ~pi221 & pi269;
assign w8821 = pi222 & ~pi270;
assign w8822 = ~w8820 & w8821;
assign w8823 = ~w8819 & ~w8822;
assign w8824 = ~w8818 & ~w8823;
assign w8825 = ~w8816 & ~w8817;
assign w8826 = ~w8824 & w8825;
assign w8827 = ~w8814 & ~w8815;
assign w8828 = ~w8826 & w8827;
assign w8829 = ~w8812 & ~w8813;
assign w8830 = ~w8828 & w8829;
assign w8831 = ~w8811 & ~w8830;
assign w8832 = ~w8810 & ~w8831;
assign w8833 = ~w8809 & ~w8832;
assign w8834 = ~w8808 & ~w8833;
assign w8835 = ~w8807 & ~w8834;
assign w8836 = ~w8806 & ~w8835;
assign w8837 = ~w8777 & w8836;
assign w8838 = pi215 & ~pi231;
assign w8839 = ~pi215 & pi231;
assign w8840 = pi216 & ~pi232;
assign w8841 = ~pi216 & pi232;
assign w8842 = pi217 & ~pi233;
assign w8843 = ~pi217 & pi233;
assign w8844 = pi218 & ~pi234;
assign w8845 = ~pi218 & pi234;
assign w8846 = pi219 & ~pi235;
assign w8847 = ~pi219 & pi235;
assign w8848 = ~pi220 & pi236;
assign w8849 = pi221 & ~pi237;
assign w8850 = ~pi221 & pi237;
assign w8851 = pi222 & ~pi238;
assign w8852 = ~w8850 & w8851;
assign w8853 = ~w8849 & ~w8852;
assign w8854 = ~w8848 & ~w8853;
assign w8855 = pi220 & ~pi236;
assign w8856 = ~w8854 & ~w8855;
assign w8857 = ~w8847 & ~w8856;
assign w8858 = ~w8846 & ~w8857;
assign w8859 = ~w8845 & ~w8858;
assign w8860 = ~w8844 & ~w8859;
assign w8861 = ~w8843 & ~w8860;
assign w8862 = ~w8842 & ~w8861;
assign w8863 = ~w8841 & ~w8862;
assign w8864 = ~w8840 & ~w8863;
assign w8865 = ~w8839 & ~w8864;
assign w8866 = ~w8838 & ~w8865;
assign w8867 = pi215 & ~pi223;
assign w8868 = ~pi215 & pi223;
assign w8869 = pi216 & ~pi224;
assign w8870 = ~pi216 & pi224;
assign w8871 = pi217 & ~pi225;
assign w8872 = ~pi217 & pi225;
assign w8873 = pi218 & ~pi226;
assign w8874 = ~pi218 & pi226;
assign w8875 = pi219 & ~pi227;
assign w8876 = ~pi219 & pi227;
assign w8877 = ~pi220 & pi228;
assign w8878 = pi221 & ~pi229;
assign w8879 = ~pi221 & pi229;
assign w8880 = pi222 & ~pi230;
assign w8881 = ~w8879 & w8880;
assign w8882 = ~w8878 & ~w8881;
assign w8883 = ~w8877 & ~w8882;
assign w8884 = pi220 & ~pi228;
assign w8885 = ~w8883 & ~w8884;
assign w8886 = ~w8876 & ~w8885;
assign w8887 = ~w8875 & ~w8886;
assign w8888 = ~w8874 & ~w8887;
assign w8889 = ~w8873 & ~w8888;
assign w8890 = ~w8872 & ~w8889;
assign w8891 = ~w8871 & ~w8890;
assign w8892 = ~w8870 & ~w8891;
assign w8893 = ~w8869 & ~w8892;
assign w8894 = ~w8868 & ~w8893;
assign w8895 = ~w8867 & ~w8894;
assign w8896 = ~pi215 & pi239;
assign w8897 = pi215 & ~pi239;
assign w8898 = ~pi216 & pi240;
assign w8899 = pi216 & ~pi240;
assign w8900 = ~pi217 & pi241;
assign w8901 = pi217 & ~pi241;
assign w8902 = pi218 & ~pi242;
assign w8903 = ~pi219 & pi243;
assign w8904 = ~pi218 & pi242;
assign w8905 = pi219 & ~pi243;
assign w8906 = pi220 & ~pi244;
assign w8907 = ~pi220 & pi244;
assign w8908 = pi221 & ~pi245;
assign w8909 = ~pi221 & pi245;
assign w8910 = pi222 & ~pi246;
assign w8911 = ~w8909 & w8910;
assign w8912 = ~w8908 & ~w8911;
assign w8913 = ~w8907 & ~w8912;
assign w8914 = ~w8905 & ~w8906;
assign w8915 = ~w8913 & w8914;
assign w8916 = ~w8903 & ~w8904;
assign w8917 = ~w8915 & w8916;
assign w8918 = ~w8901 & ~w8902;
assign w8919 = ~w8917 & w8918;
assign w8920 = ~w8900 & ~w8919;
assign w8921 = ~w8899 & ~w8920;
assign w8922 = ~w8898 & ~w8921;
assign w8923 = ~w8897 & ~w8922;
assign w8924 = ~w8896 & ~w8923;
assign w8925 = pi215 & ~pi247;
assign w8926 = ~pi215 & pi247;
assign w8927 = pi216 & ~pi248;
assign w8928 = ~pi216 & pi248;
assign w8929 = pi217 & ~pi249;
assign w8930 = ~pi218 & pi250;
assign w8931 = ~pi217 & pi249;
assign w8932 = pi218 & ~pi250;
assign w8933 = ~pi219 & pi251;
assign w8934 = pi219 & ~pi251;
assign w8935 = ~pi220 & pi252;
assign w8936 = pi220 & ~pi252;
assign w8937 = ~pi221 & pi253;
assign w8938 = pi221 & ~pi253;
assign w8939 = pi222 & ~pi254;
assign w8940 = ~w8938 & ~w8939;
assign w8941 = ~w8937 & ~w8940;
assign w8942 = ~w8936 & ~w8941;
assign w8943 = ~w8935 & ~w8942;
assign w8944 = ~w8934 & ~w8943;
assign w8945 = ~w8933 & ~w8944;
assign w8946 = ~w8932 & ~w8945;
assign w8947 = ~w8930 & ~w8931;
assign w8948 = ~w8946 & w8947;
assign w8949 = ~w8929 & ~w8948;
assign w8950 = ~w8928 & ~w8949;
assign w8951 = ~w8927 & ~w8950;
assign w8952 = ~w8926 & ~w8951;
assign w8953 = ~w8925 & ~w8952;
assign w8954 = ~w8924 & w8953;
assign w8955 = ~w206 & ~w823;
assign w8956 = w6112 & w8955;
assign w8957 = w4056 & w8001;
assign w8958 = w2594 & w7999;
assign w8959 = w8956 & w8957;
assign w8960 = w8958 & w8959;
assign w8961 = ~w1634 & w1637;
assign w8962 = w1615 & ~w8961;
assign w8963 = ~w205 & w209;
assign w8964 = ~w201 & w8963;
assign w8965 = w215 & ~w8964;
assign w8966 = w55 & w58;
assign w8967 = w33 & ~w8966;
assign w8968 = ~pi215 & ~w7000;
assign w8969 = w7997 & w8968;
assign w8970 = ~w8296 & ~w8969;
assign w8971 = ~w6070 & ~w6935;
assign w8972 = w1979 & ~w3285;
assign w8973 = w4723 & w8971;
assign w8974 = ~w8970 & w8973;
assign w8975 = ~w2071 & w8974;
assign w8976 = ~w2259 & w8960;
assign w8977 = ~w8965 & w8976;
assign w8978 = ~w8967 & w8975;
assign w8979 = w8977 & w8978;
assign w8980 = ~w1754 & ~w3165;
assign w8981 = ~w3475 & ~w4666;
assign w8982 = ~w5012 & ~w6065;
assign w8983 = ~w6929 & ~w8962;
assign w8984 = w8982 & w8983;
assign w8985 = w8980 & w8981;
assign w8986 = w8972 & w8979;
assign w8987 = w8985 & w8986;
assign w8988 = w8037 & w8984;
assign w8989 = w8987 & w8988;
assign w8990 = w8301 & w8989;
assign w8991 = w7995 & w8990;
assign w8992 = ~w7317 & w8991;
assign w8993 = w8203 & w8992;
assign w8994 = w8035 & w8837;
assign w8995 = w8866 & w8895;
assign w8996 = w8954 & w8995;
assign w8997 = w8993 & w8994;
assign w8998 = w8996 & w8997;
assign w8999 = w7647 & w17900;
assign w9000 = w5397 & w8999;
assign w9001 = pi215 & ~w6107;
assign w9002 = w2595 & ~w9001;
assign w9003 = w8748 & w9002;
assign w9004 = w8998 & w9003;
assign w9005 = w9000 & w9004;
assign w9006 = pi023 & w9005;
assign w9007 = w8342 & ~w8723;
assign w9008 = ~w8723 & w16447;
assign w9009 = (~w7648 & ~w8381) | (~w7648 & w17710) | (~w8381 & w17710);
assign w9010 = ~w6128 & w8362;
assign w9011 = ~w5738 & w9010;
assign w9012 = ~w8497 & w9011;
assign w9013 = w155 & ~w919;
assign w9014 = w597 & w2582;
assign w9015 = (w17159 & w17901) | (w17159 & w17902) | (w17901 & w17902);
assign w9016 = w9013 & w9015;
assign w9017 = w92 & w9016;
assign w9018 = w218 & w9017;
assign w9019 = ~w8659 & w9018;
assign w9020 = w8665 & w9019;
assign w9021 = w8684 & w9020;
assign w9022 = w8678 & w9021;
assign w9023 = w186 & w8347;
assign w9024 = ~w9022 & w9023;
assign w9025 = (w5432 & w7827) | (w5432 & w17903) | (w7827 & w17903);
assign w9026 = w8603 & w9025;
assign w9027 = w8618 & w9026;
assign w9028 = ~w3506 & ~w9027;
assign w9029 = ~w2902 & w8340;
assign w9030 = ~w8658 & w9029;
assign w9031 = ~w7057 & w8418;
assign w9032 = (w8031 & w16448) | (w8031 & w18478) | (w16448 & w18478);
assign w9033 = (w8294 & w16449) | (w8294 & w18478) | (w16449 & w18478);
assign w9034 = ~w9032 & w9033;
assign w9035 = ~w9031 & w9034;
assign w9036 = w7987 & w17242;
assign w9037 = w7977 & w9036;
assign w9038 = ~w9035 & ~w9037;
assign w9039 = w7198 & ~w7754;
assign w9040 = ~w4638 & w9039;
assign w9041 = (w9040 & ~w8545) | (w9040 & w16450) | (~w8545 & w16450);
assign w9042 = ~w7585 & ~w8432;
assign w9043 = ~w8432 & w16451;
assign w9044 = ~w4924 & w8344;
assign w9045 = (w9044 & ~w8492) | (w9044 & w17243) | (~w8492 & w17243);
assign w9046 = w1756 & w8653;
assign w9047 = w1727 & w8470;
assign w9048 = (w9047 & ~w8653) | (w9047 & w16452) | (~w8653 & w16452);
assign w9049 = ~w9009 & ~w9012;
assign w9050 = ~w9024 & ~w9028;
assign w9051 = ~w9030 & ~w9038;
assign w9052 = w9050 & w9051;
assign w9053 = ~w9008 & w9049;
assign w9054 = ~w9041 & ~w9043;
assign w9055 = ~w9045 & ~w9048;
assign w9056 = w9054 & w9055;
assign w9057 = w9052 & w9053;
assign w9058 = w9056 & w9057;
assign w9059 = ~pi021 & w9058;
assign w9060 = (w8368 & ~w8402) | (w8368 & w17244) | (~w8402 & w17244);
assign w9061 = w8420 & ~w8723;
assign w9062 = w8411 & ~w9022;
assign w9063 = (w8419 & ~w7977) | (w8419 & w16453) | (~w7977 & w16453);
assign w9064 = ~w3949 & ~w9027;
assign w9065 = w8416 & ~w8658;
assign w9066 = w8409 & ~w8497;
assign w9067 = (w8406 & ~w8381) | (w8406 & w17711) | (~w8381 & w17711);
assign w9068 = (w8417 & ~w8492) | (w8417 & w17245) | (~w8492 & w17245);
assign w9069 = (w7979 & ~w8333) | (w7979 & w17904) | (~w8333 & w17904);
assign w9070 = (~w7259 & ~w7992) | (~w7259 & w17905) | (~w7992 & w17905);
assign w9071 = ~w7347 & ~w8051;
assign w9072 = (w8413 & ~w8653) | (w8413 & w16454) | (~w8653 & w16454);
assign w9073 = (w8415 & ~w8545) | (w8415 & w16455) | (~w8545 & w16455);
assign w9074 = ~w5431 & w7318;
assign w9075 = w8407 & w9074;
assign w9076 = ~w9070 & w9075;
assign w9077 = ~w9071 & w9076;
assign w9078 = (w9077 & ~w8431) | (w9077 & w18341) | (~w8431 & w18341);
assign w9079 = ~w9069 & w9078;
assign w9080 = ~w9060 & ~w9061;
assign w9081 = ~w9062 & ~w9063;
assign w9082 = ~w9064 & ~w9065;
assign w9083 = ~w9066 & ~w9067;
assign w9084 = w9082 & w9083;
assign w9085 = w9080 & w9081;
assign w9086 = ~w9068 & w9079;
assign w9087 = ~w9072 & ~w9073;
assign w9088 = w9086 & w9087;
assign w9089 = w9084 & w9085;
assign w9090 = w9088 & w9089;
assign w9091 = ~pi019 & w9090;
assign w9092 = w8366 & ~w9022;
assign w9093 = w8364 & ~w8658;
assign w9094 = ~w8432 & w8369;
assign w9095 = w8365 & ~w8723;
assign w9096 = (w8367 & ~w7977) | (w8367 & w16456) | (~w7977 & w16456);
assign w9097 = w8363 & ~w8497;
assign w9098 = w3565 & ~w9027;
assign w9099 = (w8360 & ~w8492) | (w8360 & w17246) | (~w8492 & w17246);
assign w9100 = (w8370 & ~w8653) | (w8370 & w16457) | (~w8653 & w16457);
assign w9101 = (w8371 & ~w8545) | (w8371 & w16458) | (~w8545 & w16458);
assign w9102 = w9009 & ~w9060;
assign w9103 = ~w9092 & ~w9093;
assign w9104 = ~w9095 & ~w9096;
assign w9105 = ~w9097 & ~w9098;
assign w9106 = w9104 & w9105;
assign w9107 = w9102 & w9103;
assign w9108 = ~w9094 & ~w9099;
assign w9109 = ~w9100 & ~w9101;
assign w9110 = w9108 & w9109;
assign w9111 = w9106 & w9107;
assign w9112 = w9110 & w9111;
assign w9113 = w7957 & ~w8497;
assign w9114 = (w7983 & ~w8402) | (w7983 & w17247) | (~w8402 & w17247);
assign w9115 = w7978 & ~w8658;
assign w9116 = (w7980 & ~w8357) | (w7980 & w17248) | (~w8357 & w17248);
assign w9117 = (w7982 & ~w8431) | (w7982 & w17712) | (~w8431 & w17712);
assign w9118 = w7968 & ~w9022;
assign w9119 = w7962 & ~w9027;
assign w9120 = (w7964 & ~w8381) | (w7964 & w17713) | (~w8381 & w17713);
assign w9121 = w7969 & ~w8723;
assign w9122 = w8048 & w8999;
assign w9123 = w7028 & ~w9122;
assign w9124 = (w7057 & ~w7992) | (w7057 & w17906) | (~w7992 & w17906);
assign w9125 = (w7963 & ~w8545) | (w7963 & w16459) | (~w8545 & w16459);
assign w9126 = (w7970 & ~w8492) | (w7970 & w17249) | (~w8492 & w17249);
assign w9127 = (w7961 & ~w8653) | (w7961 & w16460) | (~w8653 & w16460);
assign w9128 = w7981 & ~w9124;
assign w9129 = ~w9123 & w9128;
assign w9130 = ~w7990 & w9129;
assign w9131 = ~w9113 & w9130;
assign w9132 = ~w9114 & ~w9115;
assign w9133 = ~w9116 & ~w9117;
assign w9134 = ~w9118 & ~w9119;
assign w9135 = ~w9120 & ~w9121;
assign w9136 = w9134 & w9135;
assign w9137 = w9132 & w9133;
assign w9138 = ~w9125 & w9131;
assign w9139 = ~w9126 & ~w9127;
assign w9140 = w9138 & w9139;
assign w9141 = w9136 & w9137;
assign w9142 = w9140 & w9141;
assign w9143 = ~pi017 & w9142;
assign w9144 = (w8395 & ~w8653) | (w8395 & w16461) | (~w8653 & w16461);
assign w9145 = (w8396 & ~w8545) | (w8396 & w16462) | (~w8545 & w16462);
assign w9146 = w8344 & ~w8516;
assign w9147 = (w16463 & ~w8492) | (w16463 & w17907) | (~w8492 & w17907);
assign w9148 = w8391 & ~w8497;
assign w9149 = w8393 & ~w8658;
assign w9150 = w8385 & ~w8723;
assign w9151 = w8390 & ~w9027;
assign w9152 = (w8392 & ~w7977) | (w8392 & w16464) | (~w7977 & w16464);
assign w9153 = w8394 & ~w9022;
assign w9154 = w9060 & ~w9116;
assign w9155 = ~w9148 & ~w9149;
assign w9156 = ~w9150 & ~w9151;
assign w9157 = ~w9152 & ~w9153;
assign w9158 = w9156 & w9157;
assign w9159 = w9154 & w9155;
assign w9160 = ~w9144 & ~w9145;
assign w9161 = w9159 & w9160;
assign w9162 = ~w9147 & w9158;
assign w9163 = w9161 & w9162;
assign w9164 = (w8349 & ~w8545) | (w8349 & w16465) | (~w8545 & w16465);
assign w9165 = (w8345 & ~w8492) | (w8345 & w17250) | (~w8492 & w17250);
assign w9166 = w8346 & ~w8497;
assign w9167 = w8341 & ~w8658;
assign w9168 = (w8338 & ~w8653) | (w8338 & w16466) | (~w8653 & w16466);
assign w9169 = w8343 & ~w8723;
assign w9170 = w8339 & ~w9027;
assign w9171 = ~w7967 & ~w9022;
assign w9172 = w7591 & w9171;
assign w9173 = ~w9069 & w9116;
assign w9174 = ~w9166 & ~w9167;
assign w9175 = ~w9169 & ~w9170;
assign w9176 = w9174 & w9175;
assign w9177 = ~w9164 & w9173;
assign w9178 = ~w9165 & ~w9168;
assign w9179 = ~w9172 & w9178;
assign w9180 = w9176 & w9177;
assign w9181 = w9179 & w9180;
assign w9182 = pi016 & w9181;
assign w9183 = w8340 & ~w8658;
assign w9184 = ~w8658 & w16467;
assign w9185 = w8321 & ~w9022;
assign w9186 = (w8329 & ~w8653) | (w8329 & w16468) | (~w8653 & w16468);
assign w9187 = (w8325 & ~w8545) | (w8325 & w16469) | (~w8545 & w16469);
assign w9188 = ~w3743 & ~w9027;
assign w9189 = (w8327 & ~w8492) | (w8327 & w17908) | (~w8492 & w17908);
assign w9190 = w8326 & ~w8512;
assign w9191 = w8328 & ~w8723;
assign w9192 = w9069 & ~w9190;
assign w9193 = ~w9185 & w9192;
assign w9194 = ~w9188 & ~w9191;
assign w9195 = w9193 & w9194;
assign w9196 = ~w9184 & ~w9186;
assign w9197 = ~w9187 & ~w9189;
assign w9198 = w9196 & w9197;
assign w9199 = w9195 & w9198;
assign w9200 = pi014 & w9199;
assign w9201 = w5738 & ~w8319;
assign w9202 = w5680 & ~w8051;
assign w9203 = ~w5709 & ~w9201;
assign w9204 = ~w9202 & w9203;
assign w9205 = ~w8497 & w9204;
assign w9206 = ~w9069 & w9205;
assign w9207 = ~w8723 & w16470;
assign w9208 = (w8440 & ~w8357) | (w8440 & w17251) | (~w8357 & w17251);
assign w9209 = (w8455 & ~w8545) | (w8455 & w16471) | (~w8545 & w16471);
assign w9210 = (w8443 & ~w8381) | (w8443 & w17714) | (~w8381 & w17714);
assign w9211 = w8444 & ~w9022;
assign w9212 = ~w3654 & ~w9027;
assign w9213 = w8434 & ~w8658;
assign w9214 = (w8453 & ~w8402) | (w8453 & w17909) | (~w8402 & w17909);
assign w9215 = ~w9208 & ~w9210;
assign w9216 = ~w9211 & ~w9212;
assign w9217 = ~w9213 & w9216;
assign w9218 = ~w9207 & w9215;
assign w9219 = ~w9209 & ~w9214;
assign w9220 = w9218 & w9219;
assign w9221 = w9217 & w9220;
assign w9222 = (w8470 & ~w8653) | (w8470 & w16472) | (~w8653 & w16472);
assign w9223 = ~w1329 & w9222;
assign w9224 = (w8441 & ~w8492) | (w8441 & w17252) | (~w8492 & w17252);
assign w9225 = (w8435 & ~w8431) | (w8435 & w17715) | (~w8431 & w17715);
assign w9226 = (w8454 & ~w7977) | (w8454 & w16473) | (~w7977 & w16473);
assign w9227 = ~w9225 & ~w9226;
assign w9228 = ~w9224 & w9227;
assign w9229 = ~w9223 & w9228;
assign w9230 = w8362 & w9206;
assign w9231 = w9229 & w9230;
assign w9232 = w9221 & w9231;
assign w9233 = w6376 & w9232;
assign w9234 = w6375 & ~w6416;
assign w9235 = ~w7672 & w9234;
assign w9236 = ~w9190 & w9235;
assign w9237 = w9206 & w9236;
assign w9238 = w9229 & w9237;
assign w9239 = w9221 & w9238;
assign w9240 = ~w9199 & ~w9239;
assign w9241 = w8466 & ~w9027;
assign w9242 = w8476 & ~w8658;
assign w9243 = w8478 & ~w8497;
assign w9244 = w8480 & ~w8548;
assign w9245 = ~w9241 & ~w9242;
assign w9246 = ~w9243 & w9245;
assign w9247 = ~w9244 & w9246;
assign w9248 = ~w8382 & w8475;
assign w9249 = w8477 & ~w9022;
assign w9250 = (w8472 & ~w8357) | (w8472 & w17253) | (~w8357 & w17253);
assign w9251 = ~w8403 & w8474;
assign w9252 = (w8482 & ~w7977) | (w8482 & w16474) | (~w7977 & w16474);
assign w9253 = w5377 & w9069;
assign w9254 = w4895 & ~w8051;
assign w9255 = w7992 & w8317;
assign w9256 = w4924 & ~w9255;
assign w9257 = ~w9254 & ~w9256;
assign w9258 = (w9257 & w8512) | (w9257 & w16475) | (w8512 & w16475);
assign w9259 = ~w9249 & w9258;
assign w9260 = ~w9250 & ~w9252;
assign w9261 = ~w9253 & w9260;
assign w9262 = ~w9251 & w9259;
assign w9263 = w9261 & w9262;
assign w9264 = ~w8516 & ~w9248;
assign w9265 = w9262 & w17716;
assign w9266 = (w8471 & ~w8653) | (w8471 & w16476) | (~w8653 & w16476);
assign w9267 = ~w8432 & w8465;
assign w9268 = w8481 & ~w8723;
assign w9269 = ~w9267 & ~w9268;
assign w9270 = ~w9266 & w9269;
assign w9271 = w9247 & w9270;
assign w9272 = w9265 & w9271;
assign w9273 = w8464 & w9272;
assign w9274 = ~w8497 & w8596;
assign w9275 = (w8611 & ~w7977) | (w8611 & w16477) | (~w7977 & w16477);
assign w9276 = w3534 & ~w8051;
assign w9277 = w3506 & ~w8319;
assign w9278 = ~w8512 & w8607;
assign w9279 = ~w1417 & w9222;
assign w9280 = w8606 & ~w9022;
assign w9281 = w8589 & ~w8658;
assign w9282 = ~w8432 & w8595;
assign w9283 = ~w3565 & w9009;
assign w9284 = w3478 & ~w5431;
assign w9285 = ~w9276 & w9284;
assign w9286 = ~w9277 & w9285;
assign w9287 = ~w8621 & w9286;
assign w9288 = ~w9278 & w9287;
assign w9289 = ~w9274 & ~w9275;
assign w9290 = ~w9280 & ~w9281;
assign w9291 = ~w9282 & w9290;
assign w9292 = w9288 & w9289;
assign w9293 = ~w9283 & w9292;
assign w9294 = ~w9279 & w9291;
assign w9295 = w9293 & w9294;
assign w9296 = (w8597 & ~w8492) | (w8597 & w17254) | (~w8492 & w17254);
assign w9297 = (w8604 & ~w8545) | (w8604 & w16478) | (~w8545 & w16478);
assign w9298 = (w8610 & ~w8400) | (w8610 & w17717) | (~w8400 & w17717);
assign w9299 = (w8594 & ~w8357) | (w8594 & w17256) | (~w8357 & w17256);
assign w9300 = ~w8336 & w16479;
assign w9301 = w8608 & ~w8723;
assign w9302 = ~w9298 & ~w9299;
assign w9303 = ~w9300 & ~w9301;
assign w9304 = w9302 & w9303;
assign w9305 = ~w9296 & ~w9297;
assign w9306 = w9304 & w9305;
assign w9307 = w9304 & w17718;
assign w9308 = w9295 & w9307;
assign w9309 = pi009 & w9308;
assign w9310 = w9269 & w16480;
assign w9311 = w9247 & w9310;
assign w9312 = w9265 & w9311;
assign w9313 = w8503 & ~w8548;
assign w9314 = (w8500 & ~w8653) | (w8500 & w16481) | (~w8653 & w16481);
assign w9315 = w8504 & ~w8658;
assign w9316 = (~w8499 & w8658) | (~w8499 & w16482) | (w8658 & w16482);
assign w9317 = ~w9314 & w9316;
assign w9318 = w8505 & ~w8723;
assign w9319 = w8501 & ~w9027;
assign w9320 = w8502 & ~w9022;
assign w9321 = w9190 & ~w9318;
assign w9322 = ~w9319 & ~w9320;
assign w9323 = w9321 & w9322;
assign w9324 = w9317 & w9323;
assign w9325 = w9323 & w16483;
assign w9326 = pi012 & w9325;
assign w9327 = ~w8512 & w16484;
assign w9328 = ~w8499 & ~w9327;
assign w9329 = w8524 & ~w8723;
assign w9330 = (w8529 & ~w8431) | (w8529 & w18342) | (~w8431 & w18342);
assign w9331 = ~w9329 & ~w9330;
assign w9332 = w9328 & w9331;
assign w9333 = (w8526 & ~w8492) | (w8526 & w17257) | (~w8492 & w17257);
assign w9334 = ~w8658 & w16485;
assign w9335 = (w8518 & ~w8653) | (w8518 & w16486) | (~w8653 & w16486);
assign w9336 = w8522 & ~w9027;
assign w9337 = ~w9333 & ~w9336;
assign w9338 = ~w9334 & ~w9335;
assign w9339 = w9337 & w9338;
assign w9340 = (w8527 & ~w8381) | (w8527 & w17719) | (~w8381 & w17719);
assign w9341 = w4638 & ~w8319;
assign w9342 = w4609 & ~w8051;
assign w9343 = (w8517 & ~w8357) | (w8517 & w17258) | (~w8357 & w17258);
assign w9344 = (w8528 & ~w8333) | (w8528 & w17910) | (~w8333 & w17910);
assign w9345 = (w9039 & ~w8545) | (w9039 & w16487) | (~w8545 & w16487);
assign w9346 = ~w4667 & w9345;
assign w9347 = (w8519 & ~w7977) | (w8519 & w16488) | (~w7977 & w16488);
assign w9348 = w8521 & ~w9022;
assign w9349 = ~w8497 & w8520;
assign w9350 = ~w8403 & w8530;
assign w9351 = w6519 & ~w9341;
assign w9352 = ~w9342 & w9351;
assign w9353 = ~w9344 & w9352;
assign w9354 = ~w9340 & w9353;
assign w9355 = ~w9343 & ~w9347;
assign w9356 = ~w9348 & ~w9349;
assign w9357 = ~w9350 & w9356;
assign w9358 = w9354 & w9355;
assign w9359 = w9357 & w9358;
assign w9360 = w9346 & w9359;
assign w9361 = w9331 & w16489;
assign w9362 = w9339 & w9361;
assign w9363 = w9360 & w9362;
assign w9364 = pi011 & w9363;
assign w9365 = ~w8382 & w16490;
assign w9366 = (w8570 & ~w8333) | (w8570 & w17911) | (~w8333 & w17911);
assign w9367 = w2931 & ~w8051;
assign w9368 = w2902 & ~w8319;
assign w9369 = ~w8512 & w8559;
assign w9370 = ~w8516 & w16491;
assign w9371 = w8569 & ~w9022;
assign w9372 = w8553 & ~w9027;
assign w9373 = ~w8403 & w8575;
assign w9374 = (w8573 & ~w8357) | (w8573 & w17259) | (~w8357 & w17259);
assign w9375 = (w8558 & ~w8431) | (w8558 & w17720) | (~w8431 & w17720);
assign w9376 = w8560 & ~w8723;
assign w9377 = (w8572 & ~w7977) | (w8572 & w16492) | (~w7977 & w16492);
assign w9378 = w8564 & ~w9367;
assign w9379 = ~w9368 & w9378;
assign w9380 = ~w8658 & w9379;
assign w9381 = ~w9366 & ~w9369;
assign w9382 = w9380 & w9381;
assign w9383 = ~w9371 & ~w9372;
assign w9384 = ~w9374 & ~w9375;
assign w9385 = ~w9376 & ~w9377;
assign w9386 = w9384 & w9385;
assign w9387 = w9382 & w9383;
assign w9388 = ~w9365 & ~w9373;
assign w9389 = w9387 & w9388;
assign w9390 = ~w9370 & w9386;
assign w9391 = w9389 & w9390;
assign w9392 = (w8571 & ~w8653) | (w8571 & w16493) | (~w8653 & w16493);
assign w9393 = (w8561 & ~w8545) | (w8561 & w17912) | (~w8545 & w17912);
assign w9394 = ~w8497 & w8554;
assign w9395 = ~w9392 & ~w9394;
assign w9396 = ~w9393 & w9395;
assign w9397 = w9391 & w9396;
assign w9398 = w8586 & w9397;
assign w9399 = w8552 & w9398;
assign w9400 = ~w8658 & w8712;
assign w9401 = ~w8358 & w8694;
assign w9402 = ~w8497 & w8718;
assign w9403 = ~w8432 & w8696;
assign w9404 = (w8693 & ~w8545) | (w8693 & w16494) | (~w8545 & w16494);
assign w9405 = ~w8403 & w8695;
assign w9406 = (w8691 & ~w8653) | (w8691 & w16495) | (~w8653 & w16495);
assign w9407 = ~w8516 & w8700;
assign w9408 = ~w9400 & ~w9402;
assign w9409 = ~w9405 & w9408;
assign w9410 = ~w9401 & ~w9403;
assign w9411 = ~w9404 & ~w9406;
assign w9412 = ~w9407 & w9411;
assign w9413 = w9409 & w9410;
assign w9414 = w9412 & w9413;
assign w9415 = (w8716 & ~w8381) | (w8716 & w18343) | (~w8381 & w18343);
assign w9416 = w8717 & ~w9027;
assign w9417 = w8690 & ~w9022;
assign w9418 = (w8692 & ~w7977) | (w8692 & w16496) | (~w7977 & w16496);
assign w9419 = w1981 & ~w8051;
assign w9420 = ~w7831 & ~w8699;
assign w9421 = ~w8512 & ~w9420;
assign w9422 = w2011 & ~w8319;
assign w9423 = (w8698 & ~w8333) | (w8698 & w17913) | (~w8333 & w17913);
assign w9424 = ~w4797 & ~w9419;
assign w9425 = ~w9422 & w9424;
assign w9426 = ~w8723 & w9425;
assign w9427 = ~w9421 & ~w9423;
assign w9428 = w9426 & w9427;
assign w9429 = ~w9415 & ~w9416;
assign w9430 = ~w9417 & ~w9418;
assign w9431 = w9429 & w9430;
assign w9432 = w9428 & w9431;
assign w9433 = w9431 & w16497;
assign w9434 = w9414 & w9433;
assign w9435 = pi005 & w9434;
assign w9436 = w7901 & ~w7960;
assign w9437 = w1548 & w9436;
assign w9438 = (w9437 & ~w8653) | (w9437 & w16498) | (~w8653 & w16498);
assign w9439 = w1641 & w9438;
assign w9440 = (w8634 & ~w8492) | (w8634 & w17260) | (~w8492 & w17260);
assign w9441 = ~w8497 & w9010;
assign w9442 = ~w8497 & w16499;
assign w9443 = (w8633 & ~w8545) | (w8633 & w16500) | (~w8545 & w16500);
assign w9444 = ~w9022 & w8631;
assign w9445 = ~w9440 & ~w9442;
assign w9446 = ~w9443 & ~w9444;
assign w9447 = w9445 & w9446;
assign w9448 = ~w8658 & w16501;
assign w9449 = ~w8358 & w16502;
assign w9450 = ~w8621 & w8622;
assign w9451 = ~w8512 & w16503;
assign w9452 = (w8635 & ~w7977) | (w8635 & w16504) | (~w7977 & w16504);
assign w9453 = w1137 & w9060;
assign w9454 = ~w1727 & ~w8319;
assign w9455 = (w8625 & ~w8333) | (w8625 & w17914) | (~w8333 & w17914);
assign w9456 = w1755 & ~w8051;
assign w9457 = w8628 & ~w8723;
assign w9458 = (w8630 & ~w8381) | (w8630 & w17721) | (~w8381 & w17721);
assign w9459 = ~w8432 & w8623;
assign w9460 = w7921 & ~w9454;
assign w9461 = ~w9456 & w9460;
assign w9462 = ~w9455 & w9461;
assign w9463 = ~w9450 & w9462;
assign w9464 = ~w9451 & ~w9452;
assign w9465 = ~w9457 & ~w9458;
assign w9466 = ~w9459 & w9465;
assign w9467 = w9463 & w9464;
assign w9468 = ~w9448 & ~w9449;
assign w9469 = ~w9453 & w9468;
assign w9470 = w9466 & w9467;
assign w9471 = w9469 & w9470;
assign w9472 = w1699 & w9439;
assign w9473 = w9447 & w9472;
assign w9474 = w9471 & w9473;
assign w9475 = pi003 & w9474;
assign w9476 = w7806 & w9396;
assign w9477 = w9391 & w9476;
assign w9478 = ~w186 & ~w8319;
assign w9479 = ~w217 & ~w8051;
assign w9480 = ~w4847 & ~w9478;
assign w9481 = ~w9479 & w9480;
assign w9482 = ~w9022 & w18344;
assign w9483 = ~w8516 & w16505;
assign w9484 = (w8660 & ~w8431) | (w8660 & w17722) | (~w8431 & w17722);
assign w9485 = (w8671 & ~w7977) | (w8671 & w16506) | (~w7977 & w16506);
assign w9486 = w8668 & ~w8723;
assign w9487 = ~w8621 & w8669;
assign w9488 = ~w8336 & w8672;
assign w9489 = ~w8658 & w8679;
assign w9490 = ~w8512 & w8662;
assign w9491 = (w8680 & ~w8357) | (w8680 & w17261) | (~w8357 & w17261);
assign w9492 = (w8681 & ~w8402) | (w8681 & w17262) | (~w8402 & w17262);
assign w9493 = ~w8497 & w8682;
assign w9494 = w7873 & ~w9488;
assign w9495 = ~w9490 & w9494;
assign w9496 = ~w9484 & ~w9485;
assign w9497 = ~w9486 & ~w9487;
assign w9498 = ~w9489 & ~w9491;
assign w9499 = ~w9492 & ~w9493;
assign w9500 = w9498 & w9499;
assign w9501 = w9496 & w9497;
assign w9502 = w9495 & w9501;
assign w9503 = ~w9483 & w9500;
assign w9504 = w9502 & w9503;
assign w9505 = (w8659 & ~w8381) | (w8659 & w18345) | (~w8381 & w18345);
assign w9506 = (w8670 & ~w8653) | (w8670 & w16507) | (~w8653 & w16507);
assign w9507 = (w8667 & ~w8545) | (w8667 & w17263) | (~w8545 & w17263);
assign w9508 = ~w9505 & ~w9506;
assign w9509 = ~w9507 & w9508;
assign w9510 = ~w3346 & w7184;
assign w9511 = w9482 & w9510;
assign w9512 = w9509 & w9511;
assign w9513 = w9504 & w9512;
assign w9514 = pi001 & w92;
assign w9515 = w597 & w9514;
assign w9516 = w9013 & w9515;
assign w9517 = w9513 & w9516;
assign w9518 = ~w9435 & ~w9477;
assign w9519 = ~w9475 & ~w9517;
assign w9520 = w9518 & w9519;
assign w9521 = ~w9308 & ~w9399;
assign w9522 = ~w9520 & w9521;
assign w9523 = ~w9312 & ~w9326;
assign w9524 = ~w9309 & w9523;
assign w9525 = ~w9364 & w9524;
assign w9526 = ~w9522 & w9525;
assign w9527 = w9240 & ~w9273;
assign w9528 = ~w9526 & w9527;
assign w9529 = ~w9142 & ~w9182;
assign w9530 = ~w9200 & w9529;
assign w9531 = ~w9233 & w9530;
assign w9532 = ~w9528 & w9531;
assign w9533 = ~w9143 & ~w9163;
assign w9534 = ~w9532 & w9533;
assign w9535 = pi018 & w9163;
assign w9536 = ~w9090 & ~w9535;
assign w9537 = ~w9534 & w9536;
assign w9538 = ~w9091 & ~w9112;
assign w9539 = ~w9537 & w9538;
assign w9540 = pi020 & w9112;
assign w9541 = ~w9058 & ~w9540;
assign w9542 = ~w9539 & w9541;
assign w9543 = (w8418 & ~w7977) | (w8418 & w16508) | (~w7977 & w16508);
assign w9544 = w8418 & w18479;
assign w9545 = ~w8031 & ~w8319;
assign w9546 = ~w3534 & ~w9027;
assign w9547 = w8347 & ~w9022;
assign w9548 = ~w9022 & w16509;
assign w9549 = (w7993 & ~w8431) | (w7993 & w17723) | (~w8431 & w17723);
assign w9550 = ~w8723 & w16510;
assign w9551 = ~w8497 & w16511;
assign w9552 = ~w2931 & w9183;
assign w9553 = (w16512 & ~w8492) | (w16512 & w17265) | (~w8492 & w17265);
assign w9554 = ~w4609 & w9345;
assign w9555 = ~w1755 & w9222;
assign w9556 = ~w8051 & ~w9545;
assign w9557 = (w9556 & w8382) | (w9556 & w16513) | (w8382 & w16513);
assign w9558 = ~w9546 & ~w9549;
assign w9559 = w9557 & w9558;
assign w9560 = ~w9544 & ~w9548;
assign w9561 = ~w9550 & ~w9551;
assign w9562 = ~w9552 & w9561;
assign w9563 = w9559 & w9560;
assign w9564 = ~w9553 & ~w9554;
assign w9565 = ~w9555 & w9564;
assign w9566 = w9562 & w9563;
assign w9567 = w9565 & w9566;
assign w9568 = ~w9059 & ~w9567;
assign w9569 = ~w9542 & w9568;
assign w9570 = ~w6873 & ~w7000;
assign w9571 = w8971 & w9570;
assign w9572 = w8956 & w9571;
assign w9573 = ~w957 & ~w1671;
assign w9574 = w8957 & w9573;
assign w9575 = w9572 & w9574;
assign w9576 = pi151 & w8295;
assign w9577 = ~w5014 & ~w5681;
assign w9578 = ~pi207 & w9577;
assign w9579 = ~w9576 & ~w9578;
assign w9580 = ~w2168 & ~w9579;
assign w9581 = pi223 & ~w5346;
assign w9582 = w8958 & ~w9581;
assign w9583 = ~w4059 & w5348;
assign w9584 = ~w5708 & ~w6900;
assign w9585 = ~w7565 & w9584;
assign w9586 = w7995 & w9585;
assign w9587 = w8031 & w9586;
assign w9588 = ~w7288 & w9587;
assign w9589 = ~w8291 & ~w8895;
assign w9590 = w9588 & w9589;
assign w9591 = ~w1693 & w1696;
assign w9592 = w1674 & ~w9591;
assign w9593 = ~w983 & ~w1754;
assign w9594 = ~w9592 & w9593;
assign w9595 = ~w5041 & w8033;
assign w9596 = w6103 & w9595;
assign w9597 = w2197 & ~w2259;
assign w9598 = ~w84 & w89;
assign w9599 = ~w62 & ~w9598;
assign w9600 = ~w8965 & ~w9599;
assign w9601 = ~w950 & w9600;
assign w9602 = ~w2783 & ~w3447;
assign w9603 = ~w4579 & w9602;
assign w9604 = w8972 & w9597;
assign w9605 = w9601 & w9604;
assign w9606 = w8037 & w9594;
assign w9607 = w9603 & w9606;
assign w9608 = w8301 & w9605;
assign w9609 = w9607 & w9608;
assign w9610 = w9596 & w9609;
assign w9611 = w9583 & w9610;
assign w9612 = w9590 & w9611;
assign w9613 = w4731 & w8748;
assign w9614 = w9580 & w9613;
assign w9615 = w9582 & w9614;
assign w9616 = w9575 & w9615;
assign w9617 = w9612 & w9616;
assign w9618 = ~w85 & ~w281;
assign w9619 = w4723 & w9618;
assign w9620 = w9617 & w9619;
assign w9621 = w9000 & w9620;
assign w9622 = pi024 & w9621;
assign w9623 = pi022 & w9567;
assign w9624 = ~w9006 & ~w9622;
assign w9625 = ~w9623 & w9624;
assign w9626 = ~w9569 & w9625;
assign w9627 = ~w8319 & ~w9058;
assign w9628 = ~w9058 & w16514;
assign w9629 = ~w2073 & w9007;
assign w9630 = (w9629 & ~w9414) | (w9629 & w16515) | (~w9414 & w16515);
assign w9631 = ~w9628 & ~w9630;
assign w9632 = ~w3167 & w9183;
assign w9633 = (w9632 & ~w9391) | (w9632 & w16516) | (~w9391 & w16516);
assign w9634 = (w9009 & ~w9111) | (w9009 & w17724) | (~w9111 & w17724);
assign w9635 = ~w8895 & ~w9621;
assign w9636 = w8866 & ~w9635;
assign w9637 = w8953 & ~w9005;
assign w9638 = ~w5431 & w8837;
assign w9639 = w9637 & w9638;
assign w9640 = ~w6066 & w9441;
assign w9641 = ~w9239 & w9640;
assign w9642 = ~w3477 & ~w9027;
assign w9643 = (w9642 & ~w9295) | (w9642 & w17725) | (~w9295 & w17725);
assign w9644 = ~w5013 & w9146;
assign w9645 = (w9644 & ~w9311) | (w9644 & w17726) | (~w9311 & w17726);
assign w9646 = w9017 & w9482;
assign w9647 = w9509 & w9646;
assign w9648 = w9504 & w9647;
assign w9649 = w61 & w9547;
assign w9650 = (w9649 & ~w9504) | (w9649 & w16517) | (~w9504 & w16517);
assign w9651 = ~w9641 & ~w9643;
assign w9652 = ~w9645 & ~w9650;
assign w9653 = w9651 & w9652;
assign w9654 = ~w9142 & w9543;
assign w9655 = ~w9142 & w16518;
assign w9656 = (~w9563 & w18346) | (~w9563 & w18347) | (w18346 & w18347);
assign w9657 = (w9346 & ~w9360) | (w9346 & w17727) | (~w9360 & w17727);
assign w9658 = (w9222 & ~w9471) | (w9222 & w18348) | (~w9471 & w18348);
assign w9659 = w1640 & w9658;
assign w9660 = w9042 & ~w9090;
assign w9661 = (w16520 & ~w9089) | (w16520 & w18349) | (~w9089 & w18349);
assign w9662 = ~w9655 & ~w9656;
assign w9663 = ~w9657 & ~w9661;
assign w9664 = w9662 & w9663;
assign w9665 = ~w9659 & w9664;
assign w9666 = ~w8924 & w9636;
assign w9667 = w9639 & w9666;
assign w9668 = (w9667 & w9112) | (w9667 & w16521) | (w9112 & w16521);
assign w9669 = ~w9633 & w9668;
assign w9670 = w9631 & w9669;
assign w9671 = w9653 & w9670;
assign w9672 = w9665 & w9671;
assign w9673 = (w9554 & ~w9360) | (w9554 & w17728) | (~w9360 & w17728);
assign w9674 = (w9550 & ~w9414) | (w9550 & w16522) | (~w9414 & w16522);
assign w9675 = (w9183 & ~w9391) | (w9183 & w16523) | (~w9391 & w16523);
assign w9676 = ~w2931 & w9675;
assign w9677 = (w9545 & ~w9057) | (w9545 & w17729) | (~w9057 & w17729);
assign w9678 = ~w9142 & w9544;
assign w9679 = (w9555 & ~w9471) | (w9555 & w17730) | (~w9471 & w17730);
assign w9680 = (w9549 & ~w9089) | (w9549 & w18350) | (~w9089 & w18350);
assign w9681 = (w9553 & ~w9311) | (w9553 & w17731) | (~w9311 & w17731);
assign w9682 = w9547 & ~w9648;
assign w9683 = w217 & w9682;
assign w9684 = ~w9239 & w9551;
assign w9685 = ~w9308 & w9546;
assign w9686 = ~w9634 & ~w9677;
assign w9687 = ~w9678 & ~w9680;
assign w9688 = w9686 & w9687;
assign w9689 = w9656 & ~w9673;
assign w9690 = ~w9674 & ~w9679;
assign w9691 = ~w9681 & ~w9684;
assign w9692 = ~w9685 & w9691;
assign w9693 = w9689 & w9690;
assign w9694 = ~w9676 & w9688;
assign w9695 = ~w9683 & w9694;
assign w9696 = w9692 & w9693;
assign w9697 = w9695 & w9696;
assign w9698 = ~w9672 & ~w9697;
assign w9699 = ~w8291 & ~w9621;
assign w9700 = ~w9090 & w16524;
assign w9701 = w9060 & ~w9163;
assign w9702 = w8203 & ~w9005;
assign w9703 = (w9030 & ~w9391) | (w9030 & w16525) | (~w9391 & w16525);
assign w9704 = (w9032 & ~w9566) | (w9032 & w16526) | (~w9566 & w16526);
assign w9705 = (w9045 & ~w9311) | (w9045 & w17732) | (~w9311 & w17732);
assign w9706 = (w9028 & ~w9295) | (w9028 & w17733) | (~w9295 & w17733);
assign w9707 = (w9024 & ~w9504) | (w9024 & w16527) | (~w9504 & w16527);
assign w9708 = (w9041 & ~w9360) | (w9041 & w17734) | (~w9360 & w17734);
assign w9709 = w9012 & ~w9239;
assign w9710 = (w9048 & ~w9471) | (w9048 & w17735) | (~w9471 & w17735);
assign w9711 = (w9008 & ~w9414) | (w9008 & w16528) | (~w9414 & w16528);
assign w9712 = ~w9142 & w16529;
assign w9713 = ~w9058 & w16530;
assign w9714 = w8173 & w8262;
assign w9715 = ~w9699 & w9714;
assign w9716 = ~w9702 & w9715;
assign w9717 = ~w9634 & w9716;
assign w9718 = ~w9701 & w9717;
assign w9719 = ~w9700 & ~w9703;
assign w9720 = ~w9704 & ~w9705;
assign w9721 = ~w9706 & ~w9707;
assign w9722 = ~w9708 & ~w9709;
assign w9723 = ~w9710 & ~w9711;
assign w9724 = ~w9712 & w9713;
assign w9725 = w9723 & w9724;
assign w9726 = w9721 & w9722;
assign w9727 = w9719 & w9720;
assign w9728 = w9718 & w9727;
assign w9729 = w9725 & w9726;
assign w9730 = w9728 & w9729;
assign w9731 = w9097 & ~w9239;
assign w9732 = (w9101 & ~w9360) | (w9101 & w18351) | (~w9360 & w18351);
assign w9733 = w9096 & ~w9142;
assign w9734 = (w9094 & ~w9089) | (w9094 & w18352) | (~w9089 & w18352);
assign w9735 = (w9095 & ~w9414) | (w9095 & w16531) | (~w9414 & w16531);
assign w9736 = (w9099 & ~w9311) | (w9099 & w18353) | (~w9311 & w18353);
assign w9737 = w3019 & w9675;
assign w9738 = w9098 & ~w9308;
assign w9739 = (w16532 & ~w9471) | (w16532 & w18354) | (~w9471 & w18354);
assign w9740 = (w9171 & ~w9504) | (w9171 & w16533) | (~w9504 & w16533);
assign w9741 = w9171 & w18480;
assign w9742 = w9634 & ~w9701;
assign w9743 = ~w9733 & ~w9734;
assign w9744 = w9742 & w9743;
assign w9745 = ~w9731 & ~w9732;
assign w9746 = ~w9735 & ~w9736;
assign w9747 = ~w9738 & w9746;
assign w9748 = w9744 & w9745;
assign w9749 = ~w9737 & ~w9739;
assign w9750 = ~w9741 & w9749;
assign w9751 = w9747 & w9748;
assign w9752 = w9750 & w9751;
assign w9753 = ~w9730 & ~w9752;
assign w9754 = w9698 & w9753;
assign w9755 = (w9064 & ~w9295) | (w9064 & w17736) | (~w9295 & w17736);
assign w9756 = ~w7317 & ~w9005;
assign w9757 = ~w7288 & ~w9621;
assign w9758 = (w9073 & ~w9360) | (w9073 & w17737) | (~w9360 & w17737);
assign w9759 = (w9062 & ~w9504) | (w9062 & w16534) | (~w9504 & w16534);
assign w9760 = (w9061 & ~w9414) | (w9061 & w16535) | (~w9414 & w16535);
assign w9761 = (w9072 & ~w9471) | (w9072 & w17738) | (~w9471 & w17738);
assign w9762 = w9066 & ~w9239;
assign w9763 = (w9065 & ~w9391) | (w9065 & w17739) | (~w9391 & w17739);
assign w9764 = (w9071 & ~w9566) | (w9071 & w17268) | (~w9566 & w17268);
assign w9765 = (~w8432 & ~w9089) | (~w8432 & w18355) | (~w9089 & w18355);
assign w9766 = (w9070 & ~w9057) | (w9070 & w17740) | (~w9057 & w17740);
assign w9767 = (w9068 & ~w9311) | (w9068 & w17741) | (~w9311 & w17741);
assign w9768 = w9063 & ~w9142;
assign w9769 = (w9067 & ~w9111) | (w9067 & w17742) | (~w9111 & w17742);
assign w9770 = w8407 & ~w9756;
assign w9771 = ~w9757 & w9770;
assign w9772 = (w9771 & w9163) | (w9771 & w16536) | (w9163 & w16536);
assign w9773 = w9765 & ~w9766;
assign w9774 = ~w9768 & ~w9769;
assign w9775 = w9773 & w9774;
assign w9776 = ~w9755 & w9772;
assign w9777 = ~w9758 & ~w9759;
assign w9778 = ~w9760 & ~w9761;
assign w9779 = ~w9762 & ~w9763;
assign w9780 = ~w9764 & ~w9767;
assign w9781 = w9779 & w9780;
assign w9782 = w9777 & w9778;
assign w9783 = w9775 & w9776;
assign w9784 = w9782 & w9783;
assign w9785 = w9783 & w18356;
assign w9786 = ~pi019 & w9785;
assign w9787 = (w9225 & ~w9089) | (w9225 & w18357) | (~w9089 & w18357);
assign w9788 = (w9210 & ~w9111) | (w9210 & w17743) | (~w9111 & w17743);
assign w9789 = (w9213 & ~w9391) | (w9213 & w16537) | (~w9391 & w16537);
assign w9790 = (w9212 & ~w9295) | (w9212 & w17744) | (~w9295 & w17744);
assign w9791 = (w9224 & ~w9311) | (w9224 & w17745) | (~w9311 & w17745);
assign w9792 = w9223 & ~w9474;
assign w9793 = ~w9142 & w9226;
assign w9794 = (w9201 & ~w9057) | (w9201 & w17746) | (~w9057 & w17746);
assign w9795 = ~w9163 & w9214;
assign w9796 = (w9007 & ~w9414) | (w9007 & w16538) | (~w9414 & w16538);
assign w9797 = ~w2164 & w9796;
assign w9798 = w9202 & ~w9567;
assign w9799 = w9211 & ~w9648;
assign w9800 = ~w9787 & ~w9788;
assign w9801 = ~w9793 & ~w9794;
assign w9802 = ~w9795 & w9801;
assign w9803 = ~w9789 & w9800;
assign w9804 = ~w9790 & ~w9791;
assign w9805 = ~w9792 & ~w9798;
assign w9806 = ~w9799 & w9805;
assign w9807 = w9803 & w9804;
assign w9808 = ~w9797 & w9802;
assign w9809 = w9807 & w9808;
assign w9810 = w9806 & w9809;
assign w9811 = w9209 & ~w9363;
assign w9812 = (w9116 & ~w9180) | (w9116 & w17747) | (~w9180 & w17747);
assign w9813 = w6098 & w9812;
assign w9814 = w5709 & ~w9621;
assign w9815 = w6066 & ~w9005;
assign w9816 = (w9069 & ~w9198) | (w9069 & w16539) | (~w9198 & w16539);
assign w9817 = ~w9239 & w9441;
assign w9818 = w6037 & w9817;
assign w9819 = ~w5978 & ~w9814;
assign w9820 = ~w9815 & w9819;
assign w9821 = ~w9816 & w9820;
assign w9822 = ~w9811 & w9821;
assign w9823 = ~w9813 & w9822;
assign w9824 = w9818 & w9823;
assign w9825 = w9823 & w16540;
assign w9826 = w9810 & w9825;
assign w9827 = (w9191 & ~w9414) | (w9191 & w16541) | (~w9414 & w16541);
assign w9828 = (w9184 & ~w9391) | (w9184 & w16542) | (~w9391 & w16542);
assign w9829 = (w9186 & ~w9471) | (w9186 & w17748) | (~w9471 & w17748);
assign w9830 = (w9187 & ~w9360) | (w9187 & w17749) | (~w9360 & w17749);
assign w9831 = (w9190 & ~w16483) | (w9190 & w17269) | (~w16483 & w17269);
assign w9832 = (w9189 & ~w9311) | (w9189 & w17750) | (~w9311 & w17750);
assign w9833 = (w9188 & ~w9295) | (w9188 & w17751) | (~w9295 & w17751);
assign w9834 = (w9185 & ~w9504) | (w9185 & w16543) | (~w9504 & w16543);
assign w9835 = w9816 & ~w9831;
assign w9836 = ~w9827 & w9835;
assign w9837 = ~w9828 & ~w9829;
assign w9838 = ~w9830 & ~w9832;
assign w9839 = ~w9833 & ~w9834;
assign w9840 = w9838 & w9839;
assign w9841 = w9836 & w9837;
assign w9842 = w9840 & w9841;
assign w9843 = ~w9826 & ~w9842;
assign w9844 = (w9256 & ~w9057) | (w9256 & w17752) | (~w9057 & w17752);
assign w9845 = w5013 & ~w9005;
assign w9846 = w5042 & ~w9621;
assign w9847 = (w9248 & ~w9111) | (w9248 & w17753) | (~w9111 & w17753);
assign w9848 = (w9249 & ~w9504) | (w9249 & w16544) | (~w9504 & w16544);
assign w9849 = ~w9163 & w9251;
assign w9850 = (w9250 & ~w9180) | (w9250 & w17754) | (~w9180 & w17754);
assign w9851 = ~w9142 & w9252;
assign w9852 = (w9253 & ~w9198) | (w9253 & w16545) | (~w9198 & w16545);
assign w9853 = (~w8516 & ~w9311) | (~w8516 & w17755) | (~w9311 & w17755);
assign w9854 = ~w9090 & w9267;
assign w9855 = ~w9239 & w9243;
assign w9856 = w9244 & ~w9363;
assign w9857 = w9242 & ~w9477;
assign w9858 = w9268 & ~w9434;
assign w9859 = w9254 & ~w9567;
assign w9860 = w5161 & ~w5431;
assign w9861 = ~w9845 & w9860;
assign w9862 = ~w9846 & w9861;
assign w9863 = ~w9831 & w9862;
assign w9864 = ~w9844 & ~w9847;
assign w9865 = ~w9849 & ~w9850;
assign w9866 = ~w9851 & ~w9852;
assign w9867 = w9865 & w9866;
assign w9868 = w9863 & w9864;
assign w9869 = ~w9848 & w9853;
assign w9870 = ~w9854 & ~w9855;
assign w9871 = ~w9856 & ~w9857;
assign w9872 = ~w9858 & ~w9859;
assign w9873 = w9871 & w9872;
assign w9874 = w9869 & w9870;
assign w9875 = w9867 & w9868;
assign w9876 = w9874 & w9875;
assign w9877 = w9873 & w9876;
assign w9878 = ~w1043 & w9658;
assign w9879 = w9241 & ~w9308;
assign w9880 = ~w9878 & ~w9879;
assign w9881 = w8462 & w9880;
assign w9882 = w9876 & w18358;
assign w9883 = ~pi013 & w9882;
assign w9884 = (~w9563 & w18359) | (~w9563 & w18360) | (w18359 & w18360);
assign w9885 = (w9329 & ~w9414) | (w9329 & w17270) | (~w9414 & w17270);
assign w9886 = (w9330 & ~w9089) | (w9330 & w18361) | (~w9089 & w18361);
assign w9887 = (w9348 & ~w9504) | (w9348 & w17756) | (~w9504 & w17756);
assign w9888 = w2753 & w9675;
assign w9889 = (w9333 & ~w9311) | (w9333 & w17757) | (~w9311 & w17757);
assign w9890 = ~w9474 & w17271;
assign w9891 = (w9341 & ~w9057) | (w9341 & w18362) | (~w9057 & w18362);
assign w9892 = ~w9884 & ~w9886;
assign w9893 = ~w9885 & ~w9887;
assign w9894 = ~w9889 & ~w9891;
assign w9895 = w9893 & w9894;
assign w9896 = ~w9888 & w9892;
assign w9897 = ~w9890 & w9896;
assign w9898 = w9895 & w9897;
assign w9899 = w4282 & w9345;
assign w9900 = (~w9027 & ~w9295) | (~w9027 & w18363) | (~w9295 & w18363);
assign w9901 = ~w4009 & w9900;
assign w9902 = (w9327 & ~w9323) | (w9327 & w18364) | (~w9323 & w18364);
assign w9903 = w4580 & ~w9621;
assign w9904 = w4667 & ~w9005;
assign w9905 = (w9340 & ~w9111) | (w9340 & w18365) | (~w9111 & w18365);
assign w9906 = ~w9239 & w9349;
assign w9907 = ~w9142 & w16547;
assign w9908 = (~w9198 & w17272) | (~w9198 & w17273) | (w17272 & w17273);
assign w9909 = (w9343 & ~w9180) | (w9343 & w18366) | (~w9180 & w18366);
assign w9910 = ~w9163 & w16548;
assign w9911 = w6518 & ~w8499;
assign w9912 = ~w9903 & w9911;
assign w9913 = ~w9904 & w9912;
assign w9914 = ~w9902 & w9913;
assign w9915 = ~w9363 & w9914;
assign w9916 = ~w9905 & ~w9909;
assign w9917 = w9915 & w9916;
assign w9918 = ~w9906 & ~w9907;
assign w9919 = ~w9908 & ~w9910;
assign w9920 = w9918 & w9919;
assign w9921 = w9917 & w9920;
assign w9922 = w9899 & ~w9901;
assign w9923 = w9921 & w9922;
assign w9924 = w9898 & w9923;
assign w9925 = ~pi011 & w9924;
assign w9926 = w9313 & w9324;
assign w9927 = w9363 & w9926;
assign w9928 = w9281 & ~w9477;
assign w9929 = w9280 & ~w9648;
assign w9930 = ~w9928 & ~w9929;
assign w9931 = w8592 & ~w9027;
assign w9932 = ~w9163 & w9298;
assign w9933 = w3743 & w9816;
assign w9934 = ~w9181 & w9299;
assign w9935 = ~w9112 & w9283;
assign w9936 = ~w9090 & w9282;
assign w9937 = ~w9142 & w16549;
assign w9938 = w3477 & ~w9005;
assign w9939 = w3449 & ~w9621;
assign w9940 = w3831 & ~w7757;
assign w9941 = ~w9938 & w9940;
assign w9942 = ~w9939 & w9941;
assign w9943 = (w9942 & ~w9295) | (w9942 & w17758) | (~w9295 & w17758);
assign w9944 = ~w9932 & ~w9934;
assign w9945 = ~w9936 & w9944;
assign w9946 = ~w9933 & w9943;
assign w9947 = ~w9935 & ~w9937;
assign w9948 = w9946 & w9947;
assign w9949 = w9945 & w9948;
assign w9950 = ~w9239 & w16550;
assign w9951 = (w9297 & ~w9360) | (w9297 & w17759) | (~w9360 & w17759);
assign w9952 = ~w9058 & w9277;
assign w9953 = (w9279 & ~w9471) | (w9279 & w17760) | (~w9471 & w17760);
assign w9954 = w3534 & w18481;
assign w9955 = (w9301 & ~w9414) | (w9301 & w17274) | (~w9414 & w17274);
assign w9956 = w3978 & w9831;
assign w9957 = (w9296 & ~w9311) | (w9296 & w17761) | (~w9311 & w17761);
assign w9958 = ~w9951 & ~w9952;
assign w9959 = ~w9953 & ~w9955;
assign w9960 = ~w9956 & ~w9957;
assign w9961 = w9959 & w9960;
assign w9962 = w9958 & w16551;
assign w9963 = w9961 & w9962;
assign w9964 = w9930 & w9931;
assign w9965 = w9949 & w9964;
assign w9966 = w9963 & w9965;
assign w9967 = pi009 & w9966;
assign w9968 = w7805 & w9740;
assign w9969 = w2843 & w9183;
assign w9970 = ~w3139 & ~w3254;
assign w9971 = w9969 & w9970;
assign w9972 = ~w9142 & w9377;
assign w9973 = (w9368 & ~w9057) | (w9368 & w17762) | (~w9057 & w17762);
assign w9974 = (w9375 & ~w9089) | (w9375 & w18367) | (~w9089 & w18367);
assign w9975 = (w9366 & ~w9198) | (w9366 & w16552) | (~w9198 & w16552);
assign w9976 = (w9374 & ~w9180) | (w9374 & w17763) | (~w9180 & w17763);
assign w9977 = w2784 & ~w9621;
assign w9978 = w3167 & ~w9005;
assign w9979 = ~w9163 & w9373;
assign w9980 = (w9392 & ~w9471) | (w9392 & w17764) | (~w9471 & w17764);
assign w9981 = (w9372 & ~w9295) | (w9372 & w17765) | (~w9295 & w17765);
assign w9982 = w2931 & w9656;
assign w9983 = (w16553 & ~w9111) | (w16553 & w18368) | (~w9111 & w18368);
assign w9984 = (w9376 & ~w9414) | (w9376 & w16554) | (~w9414 & w16554);
assign w9985 = (w9370 & ~w9311) | (w9370 & w17766) | (~w9311 & w17766);
assign w9986 = ~w9239 & w9394;
assign w9987 = (w9393 & ~w9360) | (w9393 & w18369) | (~w9360 & w18369);
assign w9988 = w3111 & w8562;
assign w9989 = ~w9977 & w9988;
assign w9990 = ~w9978 & w9989;
assign w9991 = ~w9369 & w9990;
assign w9992 = (w9991 & ~w9391) | (w9991 & w16555) | (~w9391 & w16555);
assign w9993 = ~w9972 & ~w9973;
assign w9994 = ~w9974 & ~w9975;
assign w9995 = ~w9976 & ~w9979;
assign w9996 = w9994 & w9995;
assign w9997 = w9992 & w9993;
assign w9998 = ~w9980 & ~w9981;
assign w9999 = ~w9983 & ~w9984;
assign w10000 = ~w9985 & ~w9986;
assign w10001 = ~w9987 & w10000;
assign w10002 = w9998 & w9999;
assign w10003 = w9996 & w9997;
assign w10004 = ~w9982 & w10003;
assign w10005 = w10001 & w10002;
assign w10006 = w10004 & w10005;
assign w10007 = (w9971 & ~w9740) | (w9971 & w18370) | (~w9740 & w18370);
assign w10008 = w10004 & w17767;
assign w10009 = (w9423 & ~w9198) | (w9423 & w16556) | (~w9198 & w16556);
assign w10010 = (w9415 & ~w9111) | (w9415 & w18371) | (~w9111 & w18371);
assign w10011 = ~w9163 & w9405;
assign w10012 = (w9403 & ~w9089) | (w9403 & w18372) | (~w9089 & w18372);
assign w10013 = ~w9142 & w9418;
assign w10014 = (w16557 & ~w9180) | (w16557 & w18373) | (~w9180 & w18373);
assign w10015 = (w9417 & ~w9504) | (w9417 & w16558) | (~w9504 & w16558);
assign w10016 = (w9406 & ~w9471) | (w9406 & w17768) | (~w9471 & w17768);
assign w10017 = ~w9239 & w9402;
assign w10018 = (w9400 & ~w9391) | (w9400 & w18374) | (~w9391 & w18374);
assign w10019 = ~w9363 & w9404;
assign w10020 = (w9198 & w9427) | (w9198 & w17275) | (w9427 & w17275);
assign w10021 = ~w10010 & ~w10011;
assign w10022 = ~w10012 & ~w10013;
assign w10023 = w10021 & w10022;
assign w10024 = ~w10014 & w10020;
assign w10025 = ~w10015 & ~w10016;
assign w10026 = ~w10017 & ~w10018;
assign w10027 = ~w10019 & w10026;
assign w10028 = w10024 & w10025;
assign w10029 = w10023 & w10028;
assign w10030 = w10027 & w10029;
assign w10031 = (w9416 & ~w9295) | (w9416 & w18375) | (~w9295 & w18375);
assign w10032 = (w9407 & ~w9311) | (w9407 & w18376) | (~w9311 & w18376);
assign w10033 = w9419 & ~w9567;
assign w10034 = w2073 & ~w9005;
assign w10035 = w2198 & ~w9621;
assign w10036 = ~w9058 & w9422;
assign w10037 = ~w4797 & ~w10034;
assign w10038 = ~w10035 & w10037;
assign w10039 = (w10038 & ~w9414) | (w10038 & w18377) | (~w9414 & w18377);
assign w10040 = ~w10036 & w10039;
assign w10041 = ~w10031 & ~w10032;
assign w10042 = ~w10033 & w10041;
assign w10043 = w10040 & w10042;
assign w10044 = w1826 & w1918;
assign w10045 = w1855 & ~w4831;
assign w10046 = ~w2103 & w10045;
assign w10047 = w6661 & w10046;
assign w10048 = w8713 & w10047;
assign w10049 = ~w8723 & w10048;
assign w10050 = w10044 & w10049;
assign w10051 = w10042 & w16559;
assign w10052 = w10030 & w10051;
assign w10053 = w1358 & w9812;
assign w10054 = (w9455 & ~w9198) | (w9455 & w17276) | (~w9198 & w17276);
assign w10055 = ~w9239 & w9442;
assign w10056 = ~w9142 & w9452;
assign w10057 = ~w10054 & ~w10056;
assign w10058 = ~w10053 & w10057;
assign w10059 = ~w10055 & w10058;
assign w10060 = (w9440 & ~w9311) | (w9440 & w17769) | (~w9311 & w17769);
assign w10061 = ~w9090 & w9459;
assign w10062 = ~w1640 & ~w9005;
assign w10063 = ~w1699 & ~w9621;
assign w10064 = w9171 & w18482;
assign w10065 = (w9450 & ~w9295) | (w9450 & w17770) | (~w9295 & w17770);
assign w10066 = (w9456 & ~w9566) | (w9456 & w16560) | (~w9566 & w16560);
assign w10067 = (w9448 & ~w9391) | (w9448 & w16561) | (~w9391 & w16561);
assign w10068 = w1168 & w9634;
assign w10069 = w7921 & ~w9474;
assign w10070 = ~w9363 & w9443;
assign w10071 = ~w9434 & w9457;
assign w10072 = (w9454 & ~w9057) | (w9454 & w17771) | (~w9057 & w17771);
assign w10073 = ~w9163 & w9453;
assign w10074 = w1611 & ~w10062;
assign w10075 = ~w10063 & w10074;
assign w10076 = ~w9451 & w10075;
assign w10077 = (w10076 & w9090) | (w10076 & w16562) | (w9090 & w16562);
assign w10078 = ~w10072 & ~w10073;
assign w10079 = w10077 & w10078;
assign w10080 = ~w10060 & ~w10065;
assign w10081 = ~w10066 & ~w10067;
assign w10082 = ~w10068 & w10069;
assign w10083 = ~w10070 & ~w10071;
assign w10084 = w10082 & w10083;
assign w10085 = w10080 & w10081;
assign w10086 = ~w10064 & w10079;
assign w10087 = w10085 & w10086;
assign w10088 = w10084 & w10087;
assign w10089 = w9438 & w10059;
assign w10090 = w10088 & w10089;
assign w10091 = w10088 & w18378;
assign w10092 = (w9479 & ~w9566) | (w9479 & w16563) | (~w9566 & w16563);
assign w10093 = (w9489 & ~w9391) | (w9489 & w16564) | (~w9391 & w16564);
assign w10094 = (w9486 & ~w9414) | (w9486 & w16565) | (~w9414 & w16565);
assign w10095 = (w9507 & ~w9360) | (w9507 & w17772) | (~w9360 & w17772);
assign w10096 = (w9487 & ~w9295) | (w9487 & w17773) | (~w9295 & w17773);
assign w10097 = ~w9239 & w9493;
assign w10098 = w852 & w9831;
assign w10099 = (w9488 & ~w9198) | (w9488 & w16566) | (~w9198 & w16566);
assign w10100 = (w9478 & ~w9057) | (w9478 & w17774) | (~w9057 & w17774);
assign w10101 = (w9506 & ~w9471) | (w9506 & w17775) | (~w9471 & w17775);
assign w10102 = ~w9112 & w9505;
assign w10103 = (w9483 & ~w9311) | (w9483 & w17776) | (~w9311 & w17776);
assign w10104 = ~w91 & ~w9621;
assign w10105 = ~w61 & ~w9005;
assign w10106 = w8661 & ~w10104;
assign w10107 = ~w10105 & w10106;
assign w10108 = (w10107 & ~w9504) | (w10107 & w16567) | (~w9504 & w16567);
assign w10109 = ~w10099 & ~w10100;
assign w10110 = ~w10102 & w10109;
assign w10111 = ~w10092 & w10108;
assign w10112 = ~w10093 & ~w10094;
assign w10113 = ~w10095 & ~w10096;
assign w10114 = ~w10097 & ~w10098;
assign w10115 = ~w10101 & ~w10103;
assign w10116 = w10114 & w10115;
assign w10117 = w10112 & w10113;
assign w10118 = w10110 & w10111;
assign w10119 = w10117 & w10118;
assign w10120 = w10116 & w10119;
assign w10121 = ~w9142 & w17278;
assign w10122 = (w9491 & ~w9180) | (w9491 & w17777) | (~w9180 & w17777);
assign w10123 = ~w9163 & w9492;
assign w10124 = ~w9090 & w9484;
assign w10125 = ~w10122 & ~w10123;
assign w10126 = ~w10124 & w10125;
assign w10127 = w9016 & ~w10121;
assign w10128 = w10126 & w10127;
assign w10129 = w9171 & w10128;
assign w10130 = w10120 & w10129;
assign w10131 = pi001 & w10130;
assign w10132 = ~w10091 & ~w10131;
assign w10133 = ~w10052 & ~w10132;
assign w10134 = pi005 & w10052;
assign w10135 = ~w10133 & ~w10134;
assign w10136 = ~w10008 & ~w10135;
assign w10137 = pi007 & w10008;
assign w10138 = ~w10136 & ~w10137;
assign w10139 = ~w9966 & ~w10138;
assign w10140 = ~w9924 & ~w9967;
assign w10141 = ~w10139 & w10140;
assign w10142 = ~w9925 & ~w9927;
assign w10143 = ~w10141 & w10142;
assign w10144 = pi012 & w9927;
assign w10145 = ~w9882 & ~w10144;
assign w10146 = ~w10143 & w10145;
assign w10147 = w9843 & ~w9883;
assign w10148 = ~w10146 & w10147;
assign w10149 = pi014 & w9842;
assign w10150 = (w9125 & ~w9360) | (w9125 & w17778) | (~w9360 & w17778);
assign w10151 = w6930 & ~w9005;
assign w10152 = w6901 & ~w9621;
assign w10153 = (w9124 & ~w9057) | (w9124 & w17779) | (~w9057 & w17779);
assign w10154 = (w9120 & ~w9111) | (w9120 & w17780) | (~w9111 & w17780);
assign w10155 = w9114 & ~w9163;
assign w10156 = (w9117 & ~w9089) | (w9117 & w18379) | (~w9089 & w18379);
assign w10157 = (w9118 & ~w9504) | (w9118 & w16568) | (~w9504 & w16568);
assign w10158 = (w9126 & ~w9311) | (w9126 & w17781) | (~w9311 & w17781);
assign w10159 = w9113 & ~w9239;
assign w10160 = (w9121 & ~w9414) | (w9121 & w16569) | (~w9414 & w16569);
assign w10161 = w6872 & ~w10151;
assign w10162 = ~w10152 & w10161;
assign w10163 = ~w7990 & w10162;
assign w10164 = (w10163 & w9181) | (w10163 & w16570) | (w9181 & w16570);
assign w10165 = ~w10153 & ~w10154;
assign w10166 = ~w10155 & ~w10156;
assign w10167 = w10165 & w10166;
assign w10168 = ~w10150 & w10164;
assign w10169 = ~w10157 & ~w10158;
assign w10170 = ~w10159 & ~w10160;
assign w10171 = w10169 & w10170;
assign w10172 = w10167 & w10168;
assign w10173 = w10171 & w10172;
assign w10174 = w6754 & w8418;
assign w10175 = ~w9142 & w10174;
assign w10176 = w6813 & w10175;
assign w10177 = (w9123 & ~w9566) | (w9123 & w16571) | (~w9566 & w16571);
assign w10178 = (w9127 & ~w9471) | (w9127 & w17782) | (~w9471 & w17782);
assign w10179 = (w9119 & ~w9295) | (w9119 & w17783) | (~w9295 & w17783);
assign w10180 = (w9115 & ~w9391) | (w9115 & w16572) | (~w9391 & w16572);
assign w10181 = ~w10177 & ~w10178;
assign w10182 = ~w10179 & ~w10180;
assign w10183 = w10181 & w10182;
assign w10184 = w10176 & w10183;
assign w10185 = w10173 & w10184;
assign w10186 = w9166 & ~w9239;
assign w10187 = (w9167 & ~w9391) | (w9167 & w16573) | (~w9391 & w16573);
assign w10188 = (w9164 & ~w9360) | (w9164 & w18380) | (~w9360 & w18380);
assign w10189 = (w9170 & ~w9295) | (w9170 & w18381) | (~w9295 & w18381);
assign w10190 = (w9168 & ~w9471) | (w9168 & w18382) | (~w9471 & w18382);
assign w10191 = (w9169 & ~w9414) | (w9169 & w16574) | (~w9414 & w16574);
assign w10192 = (w9172 & ~w9504) | (w9172 & w16575) | (~w9504 & w16575);
assign w10193 = w9812 & ~w9816;
assign w10194 = ~w10186 & w10193;
assign w10195 = ~w10187 & ~w10188;
assign w10196 = ~w10189 & ~w10190;
assign w10197 = ~w10191 & ~w10192;
assign w10198 = w10196 & w10197;
assign w10199 = w10194 & w10195;
assign w10200 = w10198 & w10199;
assign w10201 = w9146 & ~w9312;
assign w10202 = ~w5224 & w10201;
assign w10203 = w10200 & ~w10202;
assign w10204 = ~w10185 & ~w10203;
assign w10205 = pi015 & w9826;
assign w10206 = ~w10149 & w10204;
assign w10207 = ~w10205 & w10206;
assign w10208 = ~w10148 & w10207;
assign w10209 = ~pi016 & w10203;
assign w10210 = ~w9308 & w16576;
assign w10211 = w2416 & w9796;
assign w10212 = ~w9312 & w17279;
assign w10213 = (w9145 & ~w9360) | (w9145 & w17784) | (~w9360 & w17784);
assign w10214 = (w9144 & ~w9471) | (w9144 & w17785) | (~w9471 & w17785);
assign w10215 = w9148 & ~w9239;
assign w10216 = (w9149 & ~w9391) | (w9149 & w16577) | (~w9391 & w16577);
assign w10217 = ~w9142 & w9152;
assign w10218 = w9153 & ~w9648;
assign w10219 = w9701 & ~w9812;
assign w10220 = ~w10217 & w10219;
assign w10221 = ~w10213 & ~w10214;
assign w10222 = ~w10215 & ~w10216;
assign w10223 = ~w10218 & w10222;
assign w10224 = w10220 & w10221;
assign w10225 = ~w10210 & ~w10211;
assign w10226 = ~w10212 & w10225;
assign w10227 = w10223 & w10224;
assign w10228 = w10226 & w10227;
assign w10229 = ~pi017 & w10185;
assign w10230 = ~w10209 & ~w10228;
assign w10231 = ~w10229 & w10230;
assign w10232 = ~w10208 & w10231;
assign w10233 = pi018 & w10228;
assign w10234 = ~w9785 & ~w10233;
assign w10235 = ~w10232 & w10234;
assign w10236 = w9754 & ~w9786;
assign w10237 = ~w10235 & w10236;
assign w10238 = pi023 & w9672;
assign w10239 = pi021 & w9730;
assign w10240 = pi022 & w9697;
assign w10241 = pi020 & w9752;
assign w10242 = ~w10238 & ~w10239;
assign w10243 = ~w10240 & ~w10241;
assign w10244 = w10242 & w10243;
assign w10245 = ~w10237 & w10244;
assign w10246 = ~w9239 & w16578;
assign w10247 = w8895 & ~w9005;
assign w10248 = ~w9142 & w17280;
assign w10249 = ~w9058 & w17281;
assign w10250 = ~w4580 & w9345;
assign w10251 = w9332 & w9339;
assign w10252 = w9360 & w10251;
assign w10253 = (w10250 & ~w9360) | (w10250 & w18383) | (~w9360 & w18383);
assign w10254 = ~w2784 & w9675;
assign w10255 = ~w9090 & w17282;
assign w10256 = ~w2198 & w9796;
assign w10257 = (w17283 & ~w9295) | (w17283 & w18384) | (~w9295 & w18384);
assign w10258 = (w17284 & ~w9504) | (w17284 & w18385) | (~w9504 & w18385);
assign w10259 = (w17285 & ~w9311) | (w17285 & w18386) | (~w9311 & w18386);
assign w10260 = (w17286 & ~w9471) | (w17286 & w18387) | (~w9471 & w18387);
assign w10261 = ~w5431 & ~w9621;
assign w10262 = ~w10247 & w10261;
assign w10263 = (w10262 & w9163) | (w10262 & w16579) | (w9163 & w16579);
assign w10264 = ~w9656 & w10263;
assign w10265 = ~w10248 & ~w10249;
assign w10266 = ~w10253 & ~w10255;
assign w10267 = w10265 & w10266;
assign w10268 = ~w10246 & w10264;
assign w10269 = ~w10254 & ~w10256;
assign w10270 = ~w10257 & ~w10258;
assign w10271 = ~w10259 & ~w10260;
assign w10272 = w10270 & w10271;
assign w10273 = w10268 & w10269;
assign w10274 = w10267 & w10273;
assign w10275 = w10273 & w18388;
assign w10276 = ~w10245 & ~w10275;
assign w10277 = pi024 & w10275;
assign w10278 = pi231 & ~pi239;
assign w10279 = pi232 & ~pi240;
assign w10280 = ~pi232 & pi240;
assign w10281 = ~pi233 & pi241;
assign w10282 = pi233 & ~pi241;
assign w10283 = pi234 & ~pi242;
assign w10284 = ~pi234 & pi242;
assign w10285 = ~pi235 & pi243;
assign w10286 = pi235 & ~pi243;
assign w10287 = pi236 & ~pi244;
assign w10288 = ~pi237 & pi245;
assign w10289 = pi237 & ~pi245;
assign w10290 = pi238 & ~pi246;
assign w10291 = ~w10289 & ~w10290;
assign w10292 = ~pi236 & pi244;
assign w10293 = ~w10288 & ~w10292;
assign w10294 = ~w10291 & w10293;
assign w10295 = ~w10286 & ~w10287;
assign w10296 = ~w10294 & w10295;
assign w10297 = ~w10284 & ~w10285;
assign w10298 = ~w10296 & w10297;
assign w10299 = ~w10282 & ~w10283;
assign w10300 = ~w10298 & w10299;
assign w10301 = ~w10280 & ~w10281;
assign w10302 = ~w10300 & w10301;
assign w10303 = ~w10278 & ~w10279;
assign w10304 = ~w10302 & w10303;
assign w10305 = ~w111 & w115;
assign w10306 = ~w107 & w10305;
assign w10307 = w121 & ~w10306;
assign w10308 = w4712 & ~w10307;
assign w10309 = ~w10304 & w10308;
assign w10310 = w9594 & w10309;
assign w10311 = w8232 & w10310;
assign w10312 = w8924 & w10311;
assign w10313 = w7378 & w10312;
assign w10314 = w2546 & w9601;
assign w10315 = w10313 & w10314;
assign w10316 = ~w2176 & ~w9582;
assign w10317 = w8748 & ~w10316;
assign w10318 = w4730 & w10317;
assign w10319 = ~w28 & ~w2592;
assign w10320 = w9574 & w10319;
assign w10321 = ~w3081 & w9597;
assign w10322 = ~w4719 & w10321;
assign w10323 = w1609 & ~w3285;
assign w10324 = ~w4430 & w10323;
assign w10325 = ~w3799 & w10324;
assign w10326 = ~w5977 & ~w6841;
assign w10327 = w9603 & w10326;
assign w10328 = w10325 & w10327;
assign w10329 = w9590 & w10328;
assign w10330 = ~w2988 & w10329;
assign w10331 = w8038 & w10322;
assign w10332 = w10330 & w10331;
assign w10333 = ~w1790 & w1793;
assign w10334 = w1771 & ~w10333;
assign w10335 = w9583 & ~w10334;
assign w10336 = ~w5128 & w9596;
assign w10337 = ~w112 & ~w407;
assign w10338 = w9572 & w10337;
assign w10339 = w9619 & w10338;
assign w10340 = pi231 & w9576;
assign w10341 = pi239 & ~w10340;
assign w10342 = ~w2168 & ~w3055;
assign w10343 = ~w1580 & ~w1768;
assign w10344 = w10342 & w10343;
assign w10345 = ~w6814 & w9571;
assign w10346 = w10344 & w10345;
assign w10347 = ~w9579 & w10346;
assign w10348 = ~w10341 & w10347;
assign w10349 = w10320 & w10348;
assign w10350 = w10339 & w10349;
assign w10351 = w10318 & w10350;
assign w10352 = w8300 & w10351;
assign w10353 = w10336 & w10352;
assign w10354 = w10335 & w10353;
assign w10355 = w10315 & w10354;
assign w10356 = w10332 & w10355;
assign w10357 = pi026 & w10356;
assign w10358 = ~pi231 & pi247;
assign w10359 = pi231 & ~pi247;
assign w10360 = pi232 & ~pi248;
assign w10361 = ~pi233 & pi249;
assign w10362 = ~pi232 & pi248;
assign w10363 = ~pi234 & pi250;
assign w10364 = ~pi235 & pi251;
assign w10365 = pi237 & ~pi253;
assign w10366 = ~pi237 & pi253;
assign w10367 = pi238 & ~pi254;
assign w10368 = ~w10366 & w10367;
assign w10369 = ~w10365 & ~w10368;
assign w10370 = ~pi252 & ~w10369;
assign w10371 = pi235 & ~pi251;
assign w10372 = pi252 & w10369;
assign w10373 = pi236 & ~w10372;
assign w10374 = ~w10370 & ~w10371;
assign w10375 = ~w10373 & w10374;
assign w10376 = ~w10363 & ~w10364;
assign w10377 = ~w10375 & w10376;
assign w10378 = pi233 & ~pi249;
assign w10379 = pi234 & ~pi250;
assign w10380 = ~w10378 & ~w10379;
assign w10381 = ~w10377 & w10380;
assign w10382 = ~w10361 & ~w10362;
assign w10383 = ~w10381 & w10382;
assign w10384 = ~w10359 & ~w10360;
assign w10385 = ~w10383 & w10384;
assign w10386 = ~w10358 & ~w10385;
assign w10387 = ~pi231 & pi255;
assign w10388 = pi231 & ~pi255;
assign w10389 = pi232 & ~pi256;
assign w10390 = ~pi232 & pi256;
assign w10391 = ~pi233 & pi257;
assign w10392 = pi233 & ~pi257;
assign w10393 = pi234 & ~pi258;
assign w10394 = ~pi235 & pi259;
assign w10395 = ~pi234 & pi258;
assign w10396 = pi237 & ~pi261;
assign w10397 = ~pi237 & pi261;
assign w10398 = pi238 & ~pi262;
assign w10399 = ~w10397 & w10398;
assign w10400 = ~w10396 & ~w10399;
assign w10401 = ~pi260 & ~w10400;
assign w10402 = pi235 & ~pi259;
assign w10403 = pi260 & w10400;
assign w10404 = pi236 & ~w10403;
assign w10405 = ~w10401 & ~w10402;
assign w10406 = ~w10404 & w10405;
assign w10407 = ~w10394 & ~w10395;
assign w10408 = ~w10406 & w10407;
assign w10409 = ~w10392 & ~w10393;
assign w10410 = ~w10408 & w10409;
assign w10411 = ~w10390 & ~w10391;
assign w10412 = ~w10410 & w10411;
assign w10413 = ~w10388 & ~w10389;
assign w10414 = ~w10412 & w10413;
assign w10415 = ~w10387 & ~w10414;
assign w10416 = ~pi231 & pi271;
assign w10417 = pi231 & ~pi271;
assign w10418 = pi232 & ~pi272;
assign w10419 = ~pi232 & pi272;
assign w10420 = ~pi233 & pi273;
assign w10421 = pi233 & ~pi273;
assign w10422 = pi234 & ~pi274;
assign w10423 = pi235 & ~pi275;
assign w10424 = pi236 & ~pi276;
assign w10425 = ~pi237 & pi277;
assign w10426 = pi237 & ~pi277;
assign w10427 = pi238 & ~pi278;
assign w10428 = ~w10426 & ~w10427;
assign w10429 = ~pi236 & pi276;
assign w10430 = ~w10425 & ~w10429;
assign w10431 = ~w10428 & w10430;
assign w10432 = ~w10423 & ~w10424;
assign w10433 = ~w10431 & w10432;
assign w10434 = ~pi234 & pi274;
assign w10435 = ~pi235 & pi275;
assign w10436 = ~w10434 & ~w10435;
assign w10437 = ~w10433 & w10436;
assign w10438 = ~w10421 & ~w10422;
assign w10439 = ~w10437 & w10438;
assign w10440 = ~w10419 & ~w10420;
assign w10441 = ~w10439 & w10440;
assign w10442 = ~w10417 & ~w10418;
assign w10443 = ~w10441 & w10442;
assign w10444 = ~w10416 & ~w10443;
assign w10445 = ~pi231 & pi263;
assign w10446 = pi231 & ~pi263;
assign w10447 = pi232 & ~pi264;
assign w10448 = ~pi232 & pi264;
assign w10449 = ~pi233 & pi265;
assign w10450 = pi233 & ~pi265;
assign w10451 = pi234 & ~pi266;
assign w10452 = pi235 & ~pi267;
assign w10453 = pi236 & ~pi268;
assign w10454 = ~pi237 & pi269;
assign w10455 = pi237 & ~pi269;
assign w10456 = pi238 & ~pi270;
assign w10457 = ~w10455 & ~w10456;
assign w10458 = ~pi236 & pi268;
assign w10459 = ~w10454 & ~w10458;
assign w10460 = ~w10457 & w10459;
assign w10461 = ~w10452 & ~w10453;
assign w10462 = ~w10460 & w10461;
assign w10463 = ~pi234 & pi266;
assign w10464 = ~pi235 & pi267;
assign w10465 = ~w10463 & ~w10464;
assign w10466 = ~w10462 & w10465;
assign w10467 = ~w10450 & ~w10451;
assign w10468 = ~w10466 & w10467;
assign w10469 = ~w10448 & ~w10449;
assign w10470 = ~w10468 & w10469;
assign w10471 = ~w10446 & ~w10447;
assign w10472 = ~w10470 & w10471;
assign w10473 = ~w10445 & ~w10472;
assign w10474 = ~w10444 & ~w10473;
assign w10475 = ~w10386 & w10474;
assign w10476 = ~w10415 & w10475;
assign w10477 = ~pi231 & pi239;
assign w10478 = ~w10304 & ~w10477;
assign w10479 = ~w1819 & w1822;
assign w10480 = w1800 & ~w10479;
assign w10481 = ~w142 & w146;
assign w10482 = ~w138 & w10481;
assign w10483 = w152 & ~w10482;
assign w10484 = pi231 & ~w8296;
assign w10485 = w9580 & ~w10484;
assign w10486 = w1579 & w10485;
assign w10487 = ~w10483 & w10486;
assign w10488 = ~w3108 & w10487;
assign w10489 = ~w3829 & ~w5099;
assign w10490 = ~w6870 & ~w10480;
assign w10491 = w10489 & w10490;
assign w10492 = ~w10478 & w10488;
assign w10493 = w10491 & w10492;
assign w10494 = ~w4459 & ~w5946;
assign w10495 = w10493 & w10494;
assign w10496 = w10476 & w10495;
assign w10497 = ~w8261 & w10496;
assign w10498 = ~w7526 & w10497;
assign w10499 = ~w8866 & w10498;
assign w10500 = w9612 & w10499;
assign w10501 = w9575 & w10318;
assign w10502 = w10500 & w10501;
assign w10503 = ~w143 & ~w407;
assign w10504 = pi025 & w10319;
assign w10505 = w10503 & w10504;
assign w10506 = w9619 & w10505;
assign w10507 = w10502 & w10506;
assign w10508 = ~w10357 & ~w10507;
assign w10509 = w8999 & ~w10508;
assign w10510 = ~w10277 & ~w10509;
assign w10511 = ~w10276 & w10510;
assign w10512 = (w9660 & ~w9784) | (w9660 & w16580) | (~w9784 & w16580);
assign w10513 = (~w9784 & w17786) | (~w9784 & w17787) | (w17786 & w17787);
assign w10514 = w9654 & ~w10185;
assign w10515 = (w16581 & ~w10173) | (w16581 & w17788) | (~w10173 & w17788);
assign w10516 = ~w3801 & w9900;
assign w10517 = (w10516 & ~w9965) | (w10516 & w16582) | (~w9965 & w16582);
assign w10518 = w1796 & w9796;
assign w10519 = (w10518 & ~w10030) | (w10518 & w16583) | (~w10030 & w16583);
assign w10520 = w9627 & ~w9730;
assign w10521 = ~w9730 & w16584;
assign w10522 = ~w5129 & w10201;
assign w10523 = (w10522 & ~w9877) | (w10522 & w16585) | (~w9877 & w16585);
assign w10524 = ~w4431 & w9345;
assign w10525 = ~w9363 & w10524;
assign w10526 = (w10525 & ~w9923) | (w10525 & w16586) | (~w9923 & w16586);
assign w10527 = w10119 & w16587;
assign w10528 = w123 & w9682;
assign w10529 = (w10528 & ~w16587) | (w10528 & w17789) | (~w16587 & w17789);
assign w10530 = ~w3082 & w9675;
assign w10531 = (w10530 & w16588) | (w10530 & ~w10006) | (w16588 & ~w10006);
assign w10532 = w8999 & w10356;
assign w10533 = w10478 & ~w10532;
assign w10534 = ~w693 & w10320;
assign w10535 = ~w344 & w4730;
assign w10536 = w9618 & w10535;
assign w10537 = w10503 & w10536;
assign w10538 = w9572 & w10537;
assign w10539 = w10317 & w10538;
assign w10540 = w10534 & w10539;
assign w10541 = w10500 & w10540;
assign w10542 = w8999 & w10541;
assign w10543 = ~w10533 & ~w10542;
assign w10544 = ~w8924 & ~w9005;
assign w10545 = (w9658 & ~w10088) | (w9658 & w16589) | (~w10088 & w16589);
assign w10546 = (~w10088 & w17287) | (~w10088 & w17288) | (w17287 & w17288);
assign w10547 = ~w5978 & w9817;
assign w10548 = (w10547 & ~w9810) | (w10547 & w16590) | (~w9810 & w16590);
assign w10549 = (~w9621 & ~w10274) | (~w9621 & w17289) | (~w10274 & w17289);
assign w10550 = (w9656 & ~w9695) | (w9656 & w17790) | (~w9695 & w17790);
assign w10551 = (~w9748 & w18389) | (~w9748 & w18390) | (w18389 & w18390);
assign w10552 = (w9831 & ~w9363) | (w9831 & w18391) | (~w9363 & w18391);
assign w10553 = ~w8499 & ~w10552;
assign w10554 = (w9751 & w17290) | (w9751 & w17291) | (w17290 & w17291);
assign w10555 = ~w10550 & w10554;
assign w10556 = (~w10543 & w9672) | (~w10543 & w16592) | (w9672 & w16592);
assign w10557 = ~w10513 & w10556;
assign w10558 = ~w10515 & ~w10517;
assign w10559 = ~w10519 & ~w10521;
assign w10560 = ~w10523 & ~w10526;
assign w10561 = ~w10529 & ~w10531;
assign w10562 = ~w10548 & ~w10549;
assign w10563 = w10561 & w10562;
assign w10564 = w10559 & w10560;
assign w10565 = w10557 & w10558;
assign w10566 = ~w10546 & w10555;
assign w10567 = w10565 & w10566;
assign w10568 = w10563 & w10564;
assign w10569 = w10567 & w10568;
assign w10570 = (w10201 & w16593) | (w10201 & ~w9877) | (w16593 & ~w9877);
assign w10571 = ~w5100 & w10570;
assign w10572 = (w9682 & ~w16587) | (w9682 & w18392) | (~w16587 & w18392);
assign w10573 = ~w10527 & w17292;
assign w10574 = (w9796 & ~w10030) | (w9796 & w16594) | (~w10030 & w16594);
assign w10575 = w1825 & w10574;
assign w10576 = (w9900 & ~w9965) | (w9900 & w16595) | (~w9965 & w16595);
assign w10577 = ~w3830 & w10576;
assign w10578 = (w9675 & w17293) | (w9675 & ~w10006) | (w17293 & ~w10006);
assign w10579 = ~w3110 & w10578;
assign w10580 = (w9817 & ~w9810) | (w9817 & w16596) | (~w9810 & w16596);
assign w10581 = ~w5947 & w10580;
assign w10582 = ~w1579 & w10545;
assign w10583 = w7526 & w10512;
assign w10584 = (w16597 & ~w10173) | (w16597 & w18393) | (~w10173 & w18393);
assign w10585 = ~w9730 & w17294;
assign w10586 = (~w9363 & ~w9923) | (~w9363 & w16598) | (~w9923 & w16598);
assign w10587 = ~w4460 & w9345;
assign w10588 = w10586 & w10587;
assign w10589 = w8866 & ~w9005;
assign w10590 = ~w9672 & w10589;
assign w10591 = w10476 & w10543;
assign w10592 = (w10591 & w9672) | (w10591 & w16599) | (w9672 & w16599);
assign w10593 = ~w10549 & w10592;
assign w10594 = ~w10583 & ~w10584;
assign w10595 = ~w10585 & w10594;
assign w10596 = w10555 & w10593;
assign w10597 = ~w10571 & ~w10573;
assign w10598 = ~w10575 & ~w10577;
assign w10599 = ~w10579 & ~w10581;
assign w10600 = ~w10582 & ~w10588;
assign w10601 = w10599 & w10600;
assign w10602 = w10597 & w10598;
assign w10603 = w10595 & w10596;
assign w10604 = w10602 & w10603;
assign w10605 = w10601 & w10604;
assign w10606 = (w10256 & ~w10030) | (w10256 & w16600) | (~w10030 & w16600);
assign w10607 = (w10259 & w16601) | (w10259 & ~w9877) | (w16601 & ~w9877);
assign w10608 = (w10257 & ~w9965) | (w10257 & w16602) | (~w9965 & w16602);
assign w10609 = (w10260 & ~w10088) | (w10260 & w16603) | (~w10088 & w16603);
assign w10610 = (w10253 & ~w9923) | (w10253 & w16604) | (~w9923 & w16604);
assign w10611 = (w10254 & w16605) | (w10254 & ~w10006) | (w16605 & ~w10006);
assign w10612 = (w10258 & ~w16587) | (w10258 & w17791) | (~w16587 & w17791);
assign w10613 = (w10246 & ~w9810) | (w10246 & w17295) | (~w9810 & w17295);
assign w10614 = ~w9672 & w10247;
assign w10615 = ~w9730 & w10249;
assign w10616 = (w10248 & ~w10173) | (w10248 & w17792) | (~w10173 & w17792);
assign w10617 = (w10255 & ~w9784) | (w10255 & w16606) | (~w9784 & w16606);
assign w10618 = ~w10614 & ~w10615;
assign w10619 = ~w10616 & ~w10617;
assign w10620 = w10618 & w10619;
assign w10621 = w10549 & ~w10606;
assign w10622 = ~w10607 & ~w10608;
assign w10623 = ~w10609 & ~w10610;
assign w10624 = ~w10611 & ~w10612;
assign w10625 = ~w10613 & w10624;
assign w10626 = w10622 & w10623;
assign w10627 = w10620 & w16607;
assign w10628 = w10625 & w10626;
assign w10629 = w10627 & w10628;
assign w10630 = ~w10605 & ~w10629;
assign w10631 = ~w10569 & w10630;
assign w10632 = ~w6814 & w10536;
assign w10633 = w10338 & w10632;
assign w10634 = w10321 & w10633;
assign w10635 = w4722 & w10634;
assign w10636 = w10335 & w10635;
assign w10637 = w10315 & w10636;
assign w10638 = w10329 & w10637;
assign w10639 = w1915 & ~w3137;
assign w10640 = ~w4191 & w10639;
assign w10641 = ~w3771 & w10640;
assign w10642 = w8038 & w10641;
assign w10643 = w8000 & w10534;
assign w10644 = ~pi247 & pi255;
assign w10645 = pi248 & ~pi256;
assign w10646 = pi247 & ~pi255;
assign w10647 = pi249 & ~pi257;
assign w10648 = pi250 & ~pi258;
assign w10649 = ~pi250 & pi258;
assign w10650 = ~pi251 & pi259;
assign w10651 = pi251 & ~pi259;
assign w10652 = pi252 & ~pi260;
assign w10653 = ~pi253 & pi261;
assign w10654 = pi253 & ~pi261;
assign w10655 = pi254 & ~pi262;
assign w10656 = ~w10654 & ~w10655;
assign w10657 = ~pi252 & pi260;
assign w10658 = ~w10653 & ~w10657;
assign w10659 = ~w10656 & w10658;
assign w10660 = ~w10651 & ~w10652;
assign w10661 = ~w10659 & w10660;
assign w10662 = ~w10649 & ~w10650;
assign w10663 = ~w10661 & w10662;
assign w10664 = ~w10647 & ~w10648;
assign w10665 = ~w10663 & w10664;
assign w10666 = ~pi248 & pi256;
assign w10667 = ~pi249 & pi257;
assign w10668 = ~w10666 & ~w10667;
assign w10669 = ~w10665 & w10668;
assign w10670 = ~w10645 & ~w10646;
assign w10671 = ~w10669 & w10670;
assign w10672 = ~w10644 & ~w10671;
assign w10673 = pi151 & pi231;
assign w10674 = pi255 & ~w10673;
assign w10675 = w1545 & ~w5917;
assign w10676 = ~w5070 & w10675;
assign w10677 = ~w6723 & ~w10414;
assign w10678 = w10676 & w10677;
assign w10679 = w8143 & w10678;
assign w10680 = w7407 & w10679;
assign w10681 = w10336 & w10680;
assign w10682 = w8777 & w10681;
assign w10683 = pi055 & w4724;
assign w10684 = pi255 & ~w10683;
assign w10685 = ~w2756 & w10344;
assign w10686 = ~w10684 & w10685;
assign w10687 = w2549 & w2593;
assign w10688 = pi223 & ~w4714;
assign w10689 = ~w10341 & ~w10688;
assign w10690 = pi039 & pi167;
assign w10691 = w8295 & w10690;
assign w10692 = pi255 & ~w10691;
assign w10693 = ~w1729 & ~w10692;
assign w10694 = ~w530 & w10693;
assign w10695 = w10689 & w10694;
assign w10696 = w10686 & w10687;
assign w10697 = w10695 & w10696;
assign w10698 = w9577 & ~w10674;
assign w10699 = w10643 & w10698;
assign w10700 = w10672 & w10699;
assign w10701 = w10697 & w10700;
assign w10702 = w10642 & w10701;
assign w10703 = w10682 & w10702;
assign w10704 = w10638 & w10703;
assign w10705 = w8999 & w10704;
assign w10706 = pi028 & w10705;
assign w10707 = pi025 & w10605;
assign w10708 = pi024 & w10629;
assign w10709 = ~w10707 & ~w10708;
assign w10710 = ~w10569 & ~w10709;
assign w10711 = pi026 & w10569;
assign w10712 = w495 & w498;
assign w10713 = w474 & ~w10712;
assign w10714 = ~pi247 & pi271;
assign w10715 = pi247 & ~pi271;
assign w10716 = pi248 & ~pi272;
assign w10717 = pi249 & ~pi273;
assign w10718 = pi250 & ~pi274;
assign w10719 = pi251 & ~pi275;
assign w10720 = pi252 & ~pi276;
assign w10721 = ~pi253 & pi277;
assign w10722 = pi253 & ~pi277;
assign w10723 = pi254 & ~pi278;
assign w10724 = ~w10722 & ~w10723;
assign w10725 = ~pi252 & pi276;
assign w10726 = ~w10721 & ~w10725;
assign w10727 = ~w10724 & w10726;
assign w10728 = ~w10719 & ~w10720;
assign w10729 = ~w10727 & w10728;
assign w10730 = ~pi250 & pi274;
assign w10731 = ~pi251 & pi275;
assign w10732 = ~w10730 & ~w10731;
assign w10733 = ~w10729 & w10732;
assign w10734 = ~w10717 & ~w10718;
assign w10735 = ~w10733 & w10734;
assign w10736 = ~pi248 & pi272;
assign w10737 = ~pi249 & pi273;
assign w10738 = ~w10736 & ~w10737;
assign w10739 = ~w10735 & w10738;
assign w10740 = ~w10715 & ~w10716;
assign w10741 = ~w10739 & w10740;
assign w10742 = ~w10714 & ~w10741;
assign w10743 = ~pi247 & pi263;
assign w10744 = pi248 & ~pi264;
assign w10745 = pi247 & ~pi263;
assign w10746 = ~pi249 & pi265;
assign w10747 = ~pi248 & pi264;
assign w10748 = pi249 & ~pi265;
assign w10749 = pi250 & ~pi266;
assign w10750 = ~pi250 & pi266;
assign w10751 = ~pi251 & pi267;
assign w10752 = pi253 & ~pi269;
assign w10753 = ~pi253 & pi269;
assign w10754 = pi254 & ~pi270;
assign w10755 = ~w10753 & w10754;
assign w10756 = ~w10752 & ~w10755;
assign w10757 = ~pi268 & ~w10756;
assign w10758 = pi251 & ~pi267;
assign w10759 = pi268 & w10756;
assign w10760 = pi252 & ~w10759;
assign w10761 = ~w10757 & ~w10758;
assign w10762 = ~w10760 & w10761;
assign w10763 = ~w10750 & ~w10751;
assign w10764 = ~w10762 & w10763;
assign w10765 = ~w10748 & ~w10749;
assign w10766 = ~w10764 & w10765;
assign w10767 = ~w10746 & ~w10747;
assign w10768 = ~w10766 & w10767;
assign w10769 = ~w10744 & ~w10745;
assign w10770 = ~w10768 & w10769;
assign w10771 = ~w10743 & ~w10770;
assign w10772 = ~w10742 & ~w10771;
assign w10773 = ~pi247 & ~w2756;
assign w10774 = ~w5681 & w10773;
assign w10775 = ~w7108 & ~w10774;
assign w10776 = ~pi247 & ~w1580;
assign w10777 = ~w1729 & w10776;
assign w10778 = ~w6107 & ~w10777;
assign w10779 = ~w1768 & ~w5014;
assign w10780 = w10342 & w10779;
assign w10781 = w10687 & w10780;
assign w10782 = ~w10775 & w10781;
assign w10783 = ~w10778 & w10782;
assign w10784 = w1513 & w10783;
assign w10785 = w1886 & w10689;
assign w10786 = w10784 & w10785;
assign w10787 = ~w10713 & w10786;
assign w10788 = ~w4279 & ~w6035;
assign w10789 = w10643 & w10788;
assign w10790 = ~w10672 & w10787;
assign w10791 = w10789 & w10790;
assign w10792 = ~w3858 & ~w6752;
assign w10793 = w10791 & w10792;
assign w10794 = w8038 & w10386;
assign w10795 = w10793 & w10794;
assign w10796 = w8172 & w10772;
assign w10797 = w10795 & w10796;
assign w10798 = w5158 & w10336;
assign w10799 = w10797 & w10798;
assign w10800 = ~w7495 & ~w8953;
assign w10801 = w10799 & w10800;
assign w10802 = w10638 & w10801;
assign w10803 = w8999 & w10802;
assign w10804 = ~w2841 & w10803;
assign w10805 = pi027 & w10804;
assign w10806 = ~w10706 & ~w10805;
assign w10807 = ~w10711 & w10806;
assign w10808 = ~w10710 & w10807;
assign w10809 = ~w10631 & w10808;
assign w10810 = w6264 & w6271;
assign w10811 = (w16587 & w18394) | (w16587 & w18395) | (w18394 & w18395);
assign w10812 = (w9812 & ~w10200) | (w9812 & w16608) | (~w10200 & w16608);
assign w10813 = w2695 & w10812;
assign w10814 = ~w3019 & w10551;
assign w10815 = (w9984 & ~w10030) | (w9984 & w16609) | (~w10030 & w16609);
assign w10816 = ~w9697 & w9982;
assign w10817 = w3225 & w10512;
assign w10818 = ~w9730 & w9973;
assign w10819 = (w9972 & ~w10173) | (w9972 & w18396) | (~w10173 & w18396);
assign w10820 = w9968 & ~w10527;
assign w10821 = ~w10818 & ~w10819;
assign w10822 = ~w10813 & w10821;
assign w10823 = ~w10814 & ~w10815;
assign w10824 = ~w10816 & ~w10817;
assign w10825 = ~w10820 & w10824;
assign w10826 = w10822 & w10823;
assign w10827 = w10825 & w10826;
assign w10828 = w1012 & w10545;
assign w10829 = (w9978 & ~w9671) | (w9978 & w18078) | (~w9671 & w18078);
assign w10830 = w9369 & ~w9927;
assign w10831 = w3110 & ~w10542;
assign w10832 = w3082 & ~w10532;
assign w10833 = (w9979 & ~w10227) | (w9979 & w16610) | (~w10227 & w16610);
assign w10834 = w2873 & w10580;
assign w10835 = ~w9882 & w9985;
assign w10836 = ~w9966 & w9981;
assign w10837 = ~w9924 & w9987;
assign w10838 = w2784 & w10549;
assign w10839 = w8562 & ~w10831;
assign w10840 = ~w10832 & w10839;
assign w10841 = ~w9477 & w10840;
assign w10842 = ~w10830 & w10841;
assign w10843 = (w10842 & w9842) | (w10842 & w16611) | (w9842 & w16611);
assign w10844 = ~w10008 & w10843;
assign w10845 = ~w10829 & ~w10833;
assign w10846 = w10844 & w10845;
assign w10847 = ~w10835 & ~w10836;
assign w10848 = ~w10837 & w10847;
assign w10849 = ~w10828 & w10846;
assign w10850 = ~w10834 & ~w10838;
assign w10851 = w10849 & w10850;
assign w10852 = w10848 & w10851;
assign w10853 = w10826 & w16612;
assign w10854 = w10852 & w10853;
assign w10855 = ~pi007 & w10854;
assign w10856 = (w10019 & ~w9923) | (w10019 & w16613) | (~w9923 & w16613);
assign w10857 = (w10010 & ~w9751) | (w10010 & w16614) | (~w9751 & w16614);
assign w10858 = ~w9842 & w10009;
assign w10859 = ~w1825 & ~w10542;
assign w10860 = ~w1796 & ~w10532;
assign w10861 = ~w2229 & w10552;
assign w10862 = (w16615 & ~w10173) | (w16615 & w18397) | (~w10173 & w18397);
assign w10863 = (w10031 & ~w9965) | (w10031 & w16616) | (~w9965 & w16616);
assign w10864 = (~w9434 & ~w10030) | (~w9434 & w16617) | (~w10030 & w16617);
assign w10865 = (w10032 & w16618) | (w10032 & ~w9877) | (w16618 & ~w9877);
assign w10866 = (w10018 & w16619) | (w10018 & ~w10006) | (w16619 & ~w10006);
assign w10867 = w10035 & ~w10275;
assign w10868 = (~w10088 & w17297) | (~w10088 & w17298) | (w17297 & w17298);
assign w10869 = (~w9810 & w17299) | (~w9810 & w17300) | (w17299 & w17300);
assign w10870 = (w10012 & ~w9784) | (w10012 & w16620) | (~w9784 & w16620);
assign w10871 = (w10033 & ~w9695) | (w10033 & w17793) | (~w9695 & w17793);
assign w10872 = (w10036 & ~w9729) | (w10036 & w18079) | (~w9729 & w18079);
assign w10873 = (w10011 & ~w10227) | (w10011 & w16621) | (~w10227 & w16621);
assign w10874 = w7832 & ~w10859;
assign w10875 = ~w10860 & w10874;
assign w10876 = ~w10861 & w10875;
assign w10877 = ~w10858 & w10876;
assign w10878 = ~w10857 & w10877;
assign w10879 = ~w10870 & ~w10871;
assign w10880 = ~w10872 & ~w10873;
assign w10881 = w10879 & w10880;
assign w10882 = ~w10856 & w10878;
assign w10883 = ~w10862 & ~w10863;
assign w10884 = w10864 & ~w10865;
assign w10885 = ~w10866 & ~w10867;
assign w10886 = w10884 & w10885;
assign w10887 = w10882 & w10883;
assign w10888 = w10881 & w16622;
assign w10889 = w10886 & w10887;
assign w10890 = w10888 & w10889;
assign w10891 = w2444 & w10812;
assign w10892 = w9740 & ~w10527;
assign w10893 = ~w10527 & w17301;
assign w10894 = ~w9672 & w10034;
assign w10895 = ~w10891 & ~w10894;
assign w10896 = ~w10893 & w10895;
assign w10897 = w1918 & w10049;
assign w10898 = w10895 & w17302;
assign w10899 = w10889 & w16623;
assign w10900 = ~pi005 & w10899;
assign w10901 = ~w3346 & w4098;
assign w10902 = w4096 & w10901;
assign w10903 = w10120 & w16624;
assign w10904 = ~w10052 & w10094;
assign w10905 = (w10105 & ~w9671) | (w10105 & w18080) | (~w9671 & w18080);
assign w10906 = (w10124 & ~w9784) | (w10124 & w16625) | (~w9784 & w16625);
assign w10907 = w2564 & w10545;
assign w10908 = ~w9924 & w10095;
assign w10909 = (w10121 & ~w10173) | (w10121 & w17794) | (~w10173 & w17794);
assign w10910 = (w10100 & ~w9729) | (w10100 & w18081) | (~w9729 & w18081);
assign w10911 = ~w10008 & w10093;
assign w10912 = ~w913 & w10570;
assign w10913 = (w10097 & ~w9810) | (w10097 & w18398) | (~w9810 & w18398);
assign w10914 = ~w91 & w10549;
assign w10915 = ~w10905 & ~w10906;
assign w10916 = ~w10909 & ~w10910;
assign w10917 = w10915 & w10916;
assign w10918 = ~w10904 & ~w10908;
assign w10919 = ~w10911 & ~w10913;
assign w10920 = w10918 & w10919;
assign w10921 = ~w10907 & w10917;
assign w10922 = ~w10912 & ~w10914;
assign w10923 = w10921 & w10922;
assign w10924 = w10920 & w10923;
assign w10925 = w10122 & ~w10203;
assign w10926 = ~w9842 & w10099;
assign w10927 = (w10096 & ~w9965) | (w10096 & w16626) | (~w9965 & w16626);
assign w10928 = w9490 & ~w9927;
assign w10929 = (w9701 & ~w10227) | (w9701 & w16627) | (~w10227 & w16627);
assign w10930 = w659 & w10929;
assign w10931 = (w10092 & ~w9695) | (w10092 & w18399) | (~w9695 & w18399);
assign w10932 = ~w9752 & w10102;
assign w10933 = ~w123 & ~w10532;
assign w10934 = ~w154 & ~w10542;
assign w10935 = w8661 & ~w10933;
assign w10936 = ~w10934 & w10935;
assign w10937 = w9740 & w10936;
assign w10938 = ~w10928 & w10937;
assign w10939 = (w10938 & w9842) | (w10938 & w16628) | (w9842 & w16628);
assign w10940 = ~w10130 & w10939;
assign w10941 = ~w10925 & ~w10931;
assign w10942 = ~w10932 & w10941;
assign w10943 = w10940 & w16629;
assign w10944 = w10942 & w10943;
assign w10945 = w7892 & w10944;
assign w10946 = w10924 & w10945;
assign w10947 = ~w7183 & w7890;
assign w10948 = w10924 & w16630;
assign w10949 = w9451 & ~w9927;
assign w10950 = ~w9672 & w10062;
assign w10951 = ~w10008 & w10067;
assign w10952 = (w10073 & ~w10227) | (w10073 & w18400) | (~w10227 & w18400);
assign w10953 = ~w9752 & w10068;
assign w10954 = ~w9842 & w10054;
assign w10955 = w1610 & ~w10532;
assign w10956 = w1579 & ~w10542;
assign w10957 = ~w10955 & ~w10956;
assign w10958 = w10069 & w10957;
assign w10959 = ~w10954 & w10958;
assign w10960 = ~w10090 & w10959;
assign w10961 = ~w10950 & ~w10952;
assign w10962 = ~w10953 & w10961;
assign w10963 = ~w10951 & w10960;
assign w10964 = w10962 & w10963;
assign w10965 = (w10056 & ~w10173) | (w10056 & w17795) | (~w10173 & w17795);
assign w10966 = w1358 & w10812;
assign w10967 = w1329 & w10580;
assign w10968 = (w10061 & ~w9784) | (w10061 & w16631) | (~w9784 & w16631);
assign w10969 = ~w9730 & w16632;
assign w10970 = (w10060 & w16633) | (w10060 & ~w9877) | (w16633 & ~w9877);
assign w10971 = (w10064 & ~w16587) | (w10064 & w18401) | (~w16587 & w18401);
assign w10972 = w10063 & ~w10275;
assign w10973 = ~w10052 & w10071;
assign w10974 = (w10066 & ~w9695) | (w10066 & w18402) | (~w9695 & w18402);
assign w10975 = ~w9966 & w10065;
assign w10976 = ~w9924 & w10070;
assign w10977 = ~w10965 & ~w10968;
assign w10978 = ~w10974 & w10977;
assign w10979 = ~w10966 & ~w10969;
assign w10980 = ~w10970 & ~w10971;
assign w10981 = ~w10972 & ~w10973;
assign w10982 = ~w10975 & ~w10976;
assign w10983 = w10981 & w10982;
assign w10984 = w10979 & w10980;
assign w10985 = ~w10967 & w10978;
assign w10986 = w10984 & w10985;
assign w10987 = w10983 & w10986;
assign w10988 = w9438 & ~w10949;
assign w10989 = w10964 & w10988;
assign w10990 = w10987 & w10989;
assign w10991 = w10987 & w17303;
assign w10992 = ~w10899 & ~w10948;
assign w10993 = ~w10991 & w10992;
assign w10994 = ~w10900 & ~w10903;
assign w10995 = pi006 & w10903;
assign w10996 = ~w10854 & ~w10995;
assign w10997 = (w10996 & w10993) | (w10996 & w17304) | (w10993 & w17304);
assign w10998 = ~w10811 & ~w10855;
assign w10999 = ~w10997 & w10998;
assign w11000 = w9816 & ~w9842;
assign w11001 = w3743 & w11000;
assign w11002 = w3830 & ~w10542;
assign w11003 = w3801 & ~w10532;
assign w11004 = ~w3565 & w10551;
assign w11005 = w3978 & w10552;
assign w11006 = w3683 & w10812;
assign w11007 = (w9954 & ~w9695) | (w9954 & w18403) | (~w9695 & w18403);
assign w11008 = (w9932 & ~w10227) | (w9932 & w18404) | (~w10227 & w18404);
assign w11009 = (w9950 & ~w9810) | (w9950 & w16634) | (~w9810 & w16634);
assign w11010 = ~w7757 & ~w11002;
assign w11011 = ~w11003 & w11010;
assign w11012 = ~w9308 & w11011;
assign w11013 = ~w11005 & w11012;
assign w11014 = ~w9966 & w11013;
assign w11015 = ~w11001 & ~w11008;
assign w11016 = w11014 & w11015;
assign w11017 = ~w11004 & ~w11006;
assign w11018 = ~w11007 & ~w11009;
assign w11019 = w11017 & w11018;
assign w11020 = w11016 & w11019;
assign w11021 = w3714 & w10570;
assign w11022 = (w9955 & ~w10030) | (w9955 & w16635) | (~w10030 & w16635);
assign w11023 = (w9953 & ~w10088) | (w9953 & w16636) | (~w10088 & w16636);
assign w11024 = (w9952 & ~w9729) | (w9952 & w18082) | (~w9729 & w18082);
assign w11025 = (w9937 & ~w10173) | (w9937 & w17796) | (~w10173 & w17796);
assign w11026 = w9939 & ~w10275;
assign w11027 = (w9938 & ~w9671) | (w9938 & w18083) | (~w9671 & w18083);
assign w11028 = (w9936 & ~w9784) | (w9936 & w16637) | (~w9784 & w16637);
assign w11029 = w9928 & ~w10008;
assign w11030 = w9929 & ~w10527;
assign w11031 = w9297 & w10586;
assign w11032 = ~w11024 & ~w11025;
assign w11033 = ~w11027 & ~w11028;
assign w11034 = w11032 & w11033;
assign w11035 = ~w11022 & ~w11023;
assign w11036 = ~w11026 & ~w11029;
assign w11037 = ~w11030 & w11036;
assign w11038 = w11034 & w11035;
assign w11039 = ~w11021 & ~w11031;
assign w11040 = w11038 & w11039;
assign w11041 = w11037 & w11040;
assign w11042 = w11019 & w18405;
assign w11043 = w11041 & w11042;
assign w11044 = pi008 & w10811;
assign w11045 = ~w11043 & ~w11044;
assign w11046 = ~w10999 & w11045;
assign w11047 = w7785 & w7794;
assign w11048 = w10120 & w16638;
assign w11049 = ~pi009 & w11043;
assign w11050 = ~w11048 & ~w11049;
assign w11051 = ~w11046 & w11050;
assign w11052 = w9901 & ~w9966;
assign w11053 = (w9886 & ~w9784) | (w9886 & w16639) | (~w9784 & w16639);
assign w11054 = w9909 & ~w10203;
assign w11055 = ~w9672 & w9904;
assign w11056 = w4431 & ~w10532;
assign w11057 = ~w9328 & ~w10553;
assign w11058 = w4460 & ~w10542;
assign w11059 = ~w9697 & w9884;
assign w11060 = ~w11056 & ~w11058;
assign w11061 = ~w11057 & w11060;
assign w11062 = ~w11053 & w11061;
assign w11063 = ~w11054 & ~w11055;
assign w11064 = ~w11059 & w11063;
assign w11065 = w10586 & w11062;
assign w11066 = ~w11052 & w11065;
assign w11067 = w11064 & w11066;
assign w11068 = (w9910 & ~w10227) | (w9910 & w16640) | (~w10227 & w16640);
assign w11069 = (w9905 & ~w9751) | (w9905 & w16641) | (~w9751 & w16641);
assign w11070 = (w9885 & ~w10030) | (w9885 & w16642) | (~w10030 & w16642);
assign w11071 = ~w9730 & w9891;
assign w11072 = ~w9842 & w9908;
assign w11073 = (w9888 & w16643) | (w9888 & ~w10006) | (w16643 & ~w10006);
assign w11074 = (w9887 & ~w16587) | (w9887 & w18406) | (~w16587 & w18406);
assign w11075 = (w9906 & ~w9810) | (w9906 & w18407) | (~w9810 & w18407);
assign w11076 = (w9890 & ~w10088) | (w9890 & w18408) | (~w10088 & w18408);
assign w11077 = (w9907 & ~w10173) | (w9907 & w18409) | (~w10173 & w18409);
assign w11078 = ~w9882 & w9889;
assign w11079 = w4580 & w10549;
assign w11080 = ~w11068 & ~w11072;
assign w11081 = ~w11069 & ~w11071;
assign w11082 = ~w11070 & w11080;
assign w11083 = ~w11073 & ~w11074;
assign w11084 = ~w11075 & ~w11076;
assign w11085 = ~w11078 & w11084;
assign w11086 = w11082 & w11083;
assign w11087 = w11081 & w17305;
assign w11088 = w11086 & w11087;
assign w11089 = w11085 & w11088;
assign w11090 = w11066 & w18410;
assign w11091 = w11089 & w11090;
assign w11092 = pi010 & w11048;
assign w11093 = ~w11091 & ~w11092;
assign w11094 = ~w11051 & w11093;
assign w11095 = w9313 & w10586;
assign w11096 = w9318 & w10864;
assign w11097 = w9320 & ~w10527;
assign w11098 = (w9319 & ~w9965) | (w9319 & w17306) | (~w9965 & w17306);
assign w11099 = (w9317 & w10527) | (w9317 & w17307) | (w10527 & w17307);
assign w11100 = ~w11098 & w11099;
assign w11101 = ~w11095 & ~w11096;
assign w11102 = w11100 & w11101;
assign w11103 = w11101 & w17308;
assign w11104 = w6098 & w10812;
assign w11105 = (w9793 & ~w10173) | (w9793 & w18411) | (~w10173 & w18411);
assign w11106 = (w9798 & ~w9695) | (w9798 & w18412) | (~w9695 & w18412);
assign w11107 = ~w9730 & w9794;
assign w11108 = w9814 & ~w10275;
assign w11109 = (w9789 & w16644) | (w9789 & ~w10006) | (w16644 & ~w10006);
assign w11110 = (w9790 & ~w9965) | (w9790 & w16645) | (~w9965 & w16645);
assign w11111 = w9799 & ~w10527;
assign w11112 = ~w11105 & ~w11106;
assign w11113 = ~w11107 & w11112;
assign w11114 = ~w11104 & ~w11108;
assign w11115 = ~w11109 & ~w11110;
assign w11116 = ~w11111 & w11115;
assign w11117 = w11113 & w11114;
assign w11118 = w11116 & w11117;
assign w11119 = w9791 & ~w9882;
assign w11120 = w5978 & ~w10532;
assign w11121 = w5947 & ~w10542;
assign w11122 = (w10553 & w9842) | (w10553 & w16646) | (w9842 & w16646);
assign w11123 = (w9795 & ~w10227) | (w9795 & w16647) | (~w10227 & w16647);
assign w11124 = (w9815 & ~w9671) | (w9815 & w18084) | (~w9671 & w18084);
assign w11125 = (w9787 & ~w9784) | (w9787 & w16648) | (~w9784 & w16648);
assign w11126 = ~w2164 & w10574;
assign w11127 = ~w1329 & w10545;
assign w11128 = ~w5769 & w10551;
assign w11129 = w9209 & w10586;
assign w11130 = ~w5918 & ~w11120;
assign w11131 = ~w11121 & w11130;
assign w11132 = w9818 & w11131;
assign w11133 = (w11132 & ~w9810) | (w11132 & w18413) | (~w9810 & w18413);
assign w11134 = w11122 & ~w11123;
assign w11135 = ~w11124 & ~w11125;
assign w11136 = w11134 & w11135;
assign w11137 = ~w11119 & w11133;
assign w11138 = ~w11128 & w11137;
assign w11139 = ~w11126 & w11136;
assign w11140 = ~w11127 & ~w11129;
assign w11141 = w11139 & w11140;
assign w11142 = w11138 & w11141;
assign w11143 = w11117 & w16649;
assign w11144 = w11142 & w11143;
assign w11145 = (w9834 & ~w16587) | (w9834 & w17797) | (~w16587 & w17797);
assign w11146 = (w9832 & w16650) | (w9832 & ~w9877) | (w16650 & ~w9877);
assign w11147 = (w9827 & ~w10030) | (w9827 & w16651) | (~w10030 & w16651);
assign w11148 = (w9833 & ~w9965) | (w9833 & w16652) | (~w9965 & w16652);
assign w11149 = (w9829 & ~w10088) | (w9829 & w16653) | (~w10088 & w16653);
assign w11150 = (w9828 & w16654) | (w9828 & ~w10006) | (w16654 & ~w10006);
assign w11151 = (w9830 & ~w9923) | (w9830 & w16655) | (~w9923 & w16655);
assign w11152 = ~w9842 & w17309;
assign w11153 = ~w11145 & w11152;
assign w11154 = ~w11146 & ~w11147;
assign w11155 = ~w11148 & ~w11149;
assign w11156 = ~w11150 & ~w11151;
assign w11157 = w11155 & w11156;
assign w11158 = w11153 & w11154;
assign w11159 = w11157 & w11158;
assign w11160 = ~w11144 & ~w11159;
assign w11161 = (w9856 & ~w9923) | (w9856 & w16656) | (~w9923 & w16656);
assign w11162 = ~w5192 & w10512;
assign w11163 = w8466 & w10576;
assign w11164 = w9846 & ~w10275;
assign w11165 = (w16657 & ~w10173) | (w16657 & w18414) | (~w10173 & w18414);
assign w11166 = (w9878 & ~w10088) | (w9878 & w16658) | (~w10088 & w16658);
assign w11167 = (w9848 & ~w16587) | (w9848 & w18415) | (~w16587 & w18415);
assign w11168 = ~w9842 & w9852;
assign w11169 = w9850 & ~w10200;
assign w11170 = w5129 & ~w10532;
assign w11171 = w5100 & ~w10542;
assign w11172 = w9858 & ~w10052;
assign w11173 = (w9849 & ~w10227) | (w9849 & w16659) | (~w10227 & w16659);
assign w11174 = (w9844 & ~w9729) | (w9844 & w18085) | (~w9729 & w18085);
assign w11175 = (w9859 & ~w9695) | (w9859 & w17798) | (~w9695 & w17798);
assign w11176 = (w9847 & ~w9751) | (w9847 & w16660) | (~w9751 & w16660);
assign w11177 = ~w4954 & ~w5158;
assign w11178 = ~w11170 & w11177;
assign w11179 = ~w11171 & w11178;
assign w11180 = w10553 & w11179;
assign w11181 = ~w11168 & w11180;
assign w11182 = ~w11169 & w11181;
assign w11183 = ~w11173 & ~w11174;
assign w11184 = ~w11175 & ~w11176;
assign w11185 = w11183 & w11184;
assign w11186 = w10570 & w11182;
assign w11187 = ~w11161 & ~w11162;
assign w11188 = ~w11164 & ~w11165;
assign w11189 = ~w11166 & ~w11167;
assign w11190 = ~w11172 & w11189;
assign w11191 = w11187 & w11188;
assign w11192 = w11185 & w11186;
assign w11193 = ~w11163 & w11192;
assign w11194 = w11190 & w11191;
assign w11195 = w11193 & w11194;
assign w11196 = w9857 & ~w10008;
assign w11197 = ~w9826 & w9855;
assign w11198 = ~w9672 & w9845;
assign w11199 = ~w11196 & ~w11198;
assign w11200 = ~w11197 & w11199;
assign w11201 = ~w4983 & ~w5071;
assign w11202 = w11200 & w11201;
assign w11203 = w11195 & w11202;
assign w11204 = ~pi013 & w11203;
assign w11205 = w11160 & ~w11204;
assign w11206 = ~pi011 & w11091;
assign w11207 = ~w11103 & ~w11206;
assign w11208 = w11205 & w11207;
assign w11209 = ~w11094 & w11208;
assign w11210 = pi014 & w11159;
assign w11211 = pi015 & w11144;
assign w11212 = (w9769 & ~w9751) | (w9769 & w16661) | (~w9751 & w16661);
assign w11213 = (w16662 & ~w9695) | (w16662 & w18416) | (~w9695 & w18416);
assign w11214 = ~w9672 & w9756;
assign w11215 = ~w9730 & w16663;
assign w11216 = (w9768 & ~w10173) | (w9768 & w17799) | (~w10173 & w17799);
assign w11217 = ~w7526 & ~w10542;
assign w11218 = w7378 & ~w10532;
assign w11219 = (w9755 & ~w9965) | (w9755 & w16664) | (~w9965 & w16664);
assign w11220 = (w9763 & w16665) | (w9763 & ~w10006) | (w16665 & ~w10006);
assign w11221 = (w9761 & ~w10088) | (w9761 & w16666) | (~w10088 & w16666);
assign w11222 = (w9767 & w16667) | (w9767 & ~w9877) | (w16667 & ~w9877);
assign w11223 = (w9758 & ~w9923) | (w9758 & w16668) | (~w9923 & w16668);
assign w11224 = w9061 & w10864;
assign w11225 = (w10227 & w17800) | (w10227 & w17801) | (w17800 & w17801);
assign w11226 = (w9762 & ~w9810) | (w9762 & w16669) | (~w9810 & w16669);
assign w11227 = (w9759 & ~w16587) | (w9759 & w17802) | (~w16587 & w17802);
assign w11228 = w9757 & ~w10275;
assign w11229 = w7497 & ~w11217;
assign w11230 = ~w11218 & w11229;
assign w11231 = w9660 & w11230;
assign w11232 = (w11231 & ~w9784) | (w11231 & w16670) | (~w9784 & w16670);
assign w11233 = ~w11212 & w11232;
assign w11234 = ~w11214 & ~w11216;
assign w11235 = w11233 & w11234;
assign w11236 = ~w11213 & ~w11215;
assign w11237 = ~w11219 & ~w11220;
assign w11238 = ~w11221 & ~w11222;
assign w11239 = ~w11223 & w11225;
assign w11240 = ~w11226 & w18417;
assign w11241 = w11238 & w11239;
assign w11242 = w11236 & w11237;
assign w11243 = ~w11224 & w11235;
assign w11244 = w11242 & w11243;
assign w11245 = w11240 & w11241;
assign w11246 = w11244 & w11245;
assign w11247 = ~w5857 & w10580;
assign w11248 = (w10211 & ~w10030) | (w10211 & w16671) | (~w10030 & w16671);
assign w11249 = (w10216 & w16672) | (w10216 & ~w10006) | (w16672 & ~w10006);
assign w11250 = (w10218 & ~w16587) | (w10218 & w18418) | (~w16587 & w18418);
assign w11251 = (w10213 & ~w9923) | (w10213 & w16673) | (~w9923 & w16673);
assign w11252 = (w10212 & w16674) | (w10212 & ~w9877) | (w16674 & ~w9877);
assign w11253 = (w10200 & w17310) | (w10200 & w17311) | (w17310 & w17311);
assign w11254 = (w10214 & ~w10088) | (w10214 & w18419) | (~w10088 & w18419);
assign w11255 = (w10217 & ~w10173) | (w10217 & w17803) | (~w10173 & w17803);
assign w11256 = ~w9966 & w10210;
assign w11257 = w10929 & ~w11255;
assign w11258 = ~w11248 & w11257;
assign w11259 = ~w11249 & ~w11250;
assign w11260 = ~w11251 & ~w11252;
assign w11261 = w11253 & ~w11254;
assign w11262 = ~w11256 & w11261;
assign w11263 = w11259 & w11260;
assign w11264 = ~w11247 & w11258;
assign w11265 = w11263 & w11264;
assign w11266 = w11262 & w11265;
assign w11267 = ~w11246 & ~w11266;
assign w11268 = ~pi018 & ~w11246;
assign w11269 = ~w11267 & ~w11268;
assign w11270 = ~w9672 & w10151;
assign w11271 = ~w5799 & w10580;
assign w11272 = w11253 & ~w11270;
assign w11273 = ~w11271 & w11272;
assign w11274 = (w10160 & ~w10030) | (w10160 & w16675) | (~w10030 & w16675);
assign w11275 = (w10180 & w16676) | (w10180 & ~w10006) | (w16676 & ~w10006);
assign w11276 = (w16598 & w17804) | (w16598 & w17805) | (w17804 & w17805);
assign w11277 = (w10177 & ~w9695) | (w10177 & w17806) | (~w9695 & w17806);
assign w11278 = (w10153 & ~w9729) | (w10153 & w18086) | (~w9729 & w18086);
assign w11279 = (w10179 & ~w9965) | (w10179 & w16677) | (~w9965 & w16677);
assign w11280 = (w10155 & ~w10227) | (w10155 & w16678) | (~w10227 & w16678);
assign w11281 = (w10156 & ~w9784) | (w10156 & w16679) | (~w9784 & w16679);
assign w11282 = w6901 & w10549;
assign w11283 = (w10154 & ~w9751) | (w10154 & w16680) | (~w9751 & w16680);
assign w11284 = w6871 & ~w10542;
assign w11285 = w6842 & ~w10532;
assign w11286 = (w10158 & w16681) | (w10158 & ~w9877) | (w16681 & ~w9877);
assign w11287 = (w10178 & ~w10088) | (w10178 & w16682) | (~w10088 & w16682);
assign w11288 = w10157 & ~w10527;
assign w11289 = ~w5431 & ~w11284;
assign w11290 = ~w11285 & w11289;
assign w11291 = ~w7990 & w11290;
assign w11292 = (w11291 & ~w10173) | (w11291 & w17807) | (~w10173 & w17807);
assign w11293 = ~w11277 & w11292;
assign w11294 = ~w11278 & ~w11280;
assign w11295 = ~w11281 & ~w11283;
assign w11296 = w11294 & w11295;
assign w11297 = ~w11274 & w11293;
assign w11298 = ~w11275 & ~w11279;
assign w11299 = ~w11286 & ~w11287;
assign w11300 = ~w11288 & w11299;
assign w11301 = w11297 & w11298;
assign w11302 = w11296 & w16683;
assign w11303 = w11300 & w11301;
assign w11304 = w11302 & w11303;
assign w11305 = w11272 & w17314;
assign w11306 = w11303 & w16684;
assign w11307 = (w10202 & ~w9877) | (w10202 & w16685) | (~w9877 & w16685);
assign w11308 = (w10192 & ~w16587) | (w10192 & w18420) | (~w16587 & w18420);
assign w11309 = (w10191 & ~w10030) | (w10191 & w16686) | (~w10030 & w16686);
assign w11310 = (w10190 & ~w10088) | (w10190 & w17315) | (~w10088 & w17315);
assign w11311 = (w10187 & ~w10006) | (w10187 & w17316) | (~w10006 & w17316);
assign w11312 = ~w9924 & w10188;
assign w11313 = ~w6098 & w10580;
assign w11314 = ~w3683 & w10576;
assign w11315 = w10812 & w11122;
assign w11316 = ~w11307 & w11315;
assign w11317 = ~w11308 & ~w11309;
assign w11318 = ~w11310 & ~w11311;
assign w11319 = ~w11312 & w11318;
assign w11320 = w11316 & w11317;
assign w11321 = ~w11313 & ~w11314;
assign w11322 = w11320 & w11321;
assign w11323 = w11319 & w11322;
assign w11324 = ~w11306 & ~w11323;
assign w11325 = ~pi012 & ~w11203;
assign w11326 = ~w11103 & ~w11203;
assign w11327 = ~w11325 & ~w11326;
assign w11328 = w11205 & w11327;
assign w11329 = ~w11210 & ~w11211;
assign w11330 = ~w11269 & w11324;
assign w11331 = w11329 & w11330;
assign w11332 = ~w11328 & w11331;
assign w11333 = ~w11209 & w11332;
assign w11334 = (w9709 & ~w9810) | (w9709 & w16687) | (~w9810 & w16687);
assign w11335 = (w9704 & ~w9695) | (w9704 & w17808) | (~w9695 & w17808);
assign w11336 = (w9706 & ~w9965) | (w9706 & w16688) | (~w9965 & w16688);
assign w11337 = (w9707 & ~w16587) | (w9707 & w17809) | (~w16587 & w17809);
assign w11338 = (w9699 & ~w10274) | (w9699 & w17317) | (~w10274 & w17317);
assign w11339 = (w9708 & ~w9923) | (w9708 & w16689) | (~w9923 & w16689);
assign w11340 = (~w10004 & w17810) | (~w10004 & w17811) | (w17810 & w17811);
assign w11341 = (w9711 & ~w10030) | (w9711 & w16691) | (~w10030 & w16691);
assign w11342 = ~w8261 & ~w10542;
assign w11343 = w8232 & ~w10532;
assign w11344 = ~w4924 & w10570;
assign w11345 = w1727 & w10545;
assign w11346 = (w9712 & ~w10173) | (w9712 & w17812) | (~w10173 & w17812);
assign w11347 = (w9702 & ~w9671) | (w9702 & w18087) | (~w9671 & w18087);
assign w11348 = w9700 & ~w9785;
assign w11349 = w8174 & ~w11342;
assign w11350 = ~w11343 & w11349;
assign w11351 = ~w9730 & w16692;
assign w11352 = ~w10929 & ~w11335;
assign w11353 = ~w11346 & ~w11347;
assign w11354 = ~w11348 & w11353;
assign w11355 = w11351 & w11352;
assign w11356 = w10554 & ~w11334;
assign w11357 = ~w11336 & ~w11337;
assign w11358 = ~w11338 & ~w11339;
assign w11359 = ~w11340 & ~w11341;
assign w11360 = w11358 & w11359;
assign w11361 = w11356 & w11357;
assign w11362 = w11354 & w11355;
assign w11363 = ~w11344 & ~w11345;
assign w11364 = w11362 & w11363;
assign w11365 = w11360 & w11361;
assign w11366 = w11364 & w11365;
assign w11367 = (w9737 & w16693) | (w9737 & ~w10006) | (w16693 & ~w10006);
assign w11368 = (w9732 & ~w9923) | (w9732 & w16694) | (~w9923 & w16694);
assign w11369 = w3565 & w10576;
assign w11370 = (w9735 & ~w10030) | (w9735 & w16695) | (~w10030 & w16695);
assign w11371 = (w9736 & w16696) | (w9736 & ~w9877) | (w16696 & ~w9877);
assign w11372 = (w9739 & ~w10088) | (w9739 & w16697) | (~w10088 & w16697);
assign w11373 = w249 & w10572;
assign w11374 = w5769 & w10580;
assign w11375 = (w9733 & ~w10173) | (w9733 & w17813) | (~w10173 & w17813);
assign w11376 = w9734 & ~w9785;
assign w11377 = w10551 & ~w11375;
assign w11378 = ~w11376 & w11377;
assign w11379 = w11225 & ~w11367;
assign w11380 = ~w11368 & ~w11370;
assign w11381 = ~w11371 & ~w11372;
assign w11382 = w11380 & w11381;
assign w11383 = w11378 & w11379;
assign w11384 = ~w11369 & ~w11373;
assign w11385 = ~w11374 & w11384;
assign w11386 = w11382 & w11383;
assign w11387 = w11385 & w11386;
assign w11388 = ~w11366 & ~w11387;
assign w11389 = (w9676 & ~w10006) | (w9676 & w16698) | (~w10006 & w16698);
assign w11390 = w9677 & ~w9730;
assign w11391 = (w9680 & ~w9784) | (w9680 & w16699) | (~w9784 & w16699);
assign w11392 = (w9678 & ~w10173) | (w9678 & w17814) | (~w10173 & w17814);
assign w11393 = (w9674 & ~w10030) | (w9674 & w16700) | (~w10030 & w16700);
assign w11394 = (w9681 & ~w9877) | (w9681 & w16701) | (~w9877 & w16701);
assign w11395 = (w9673 & ~w9923) | (w9673 & w16702) | (~w9923 & w16702);
assign w11396 = w9683 & ~w10527;
assign w11397 = w9679 & ~w10090;
assign w11398 = w9685 & ~w9966;
assign w11399 = w9684 & ~w9826;
assign w11400 = w10550 & ~w11390;
assign w11401 = ~w11391 & ~w11392;
assign w11402 = w11400 & w11401;
assign w11403 = w10554 & ~w11389;
assign w11404 = ~w11393 & ~w11394;
assign w11405 = ~w11395 & ~w11396;
assign w11406 = ~w11397 & ~w11398;
assign w11407 = ~w11399 & w11406;
assign w11408 = w11404 & w11405;
assign w11409 = w11402 & w11403;
assign w11410 = w11408 & w11409;
assign w11411 = w11407 & w11410;
assign w11412 = (w9641 & ~w9810) | (w9641 & w16703) | (~w9810 & w16703);
assign w11413 = (w9650 & ~w10120) | (w9650 & w16704) | (~w10120 & w16704);
assign w11414 = (w9659 & ~w10088) | (w9659 & w16705) | (~w10088 & w16705);
assign w11415 = (w9657 & ~w9923) | (w9657 & w16706) | (~w9923 & w16706);
assign w11416 = (w9635 & ~w10274) | (w9635 & w17318) | (~w10274 & w17318);
assign w11417 = (w9643 & ~w9965) | (w9643 & w16707) | (~w9965 & w16707);
assign w11418 = (w9633 & w16708) | (w9633 & ~w10006) | (w16708 & ~w10006);
assign w11419 = (w9645 & w16709) | (w9645 & ~w9877) | (w16709 & ~w9877);
assign w11420 = (w9630 & ~w10030) | (w9630 & w17319) | (~w10030 & w17319);
assign w11421 = (w9628 & ~w9729) | (w9628 & w18088) | (~w9729 & w18088);
assign w11422 = ~w8866 & ~w10542;
assign w11423 = w8924 & ~w10532;
assign w11424 = (w9661 & ~w9784) | (w9661 & w16710) | (~w9784 & w16710);
assign w11425 = (w9655 & ~w10173) | (w9655 & w17815) | (~w10173 & w17815);
assign w11426 = ~w11422 & ~w11423;
assign w11427 = w9639 & w11426;
assign w11428 = (w11427 & ~w9671) | (w11427 & w18089) | (~w9671 & w18089);
assign w11429 = ~w11421 & w11428;
assign w11430 = ~w11424 & ~w11425;
assign w11431 = w11429 & w11430;
assign w11432 = ~w11412 & ~w11413;
assign w11433 = ~w11414 & ~w11415;
assign w11434 = ~w11416 & ~w11417;
assign w11435 = ~w11418 & ~w11419;
assign w11436 = ~w11420 & w11435;
assign w11437 = w11433 & w11434;
assign w11438 = w11431 & w16711;
assign w11439 = w11436 & w11437;
assign w11440 = w11438 & w11439;
assign w11441 = ~w11411 & ~w11440;
assign w11442 = w11388 & w11441;
assign w11443 = pi017 & w11306;
assign w11444 = pi016 & ~w11306;
assign w11445 = ~w11324 & ~w11443;
assign w11446 = ~w11444 & w11445;
assign w11447 = ~w11266 & ~w11446;
assign w11448 = ~w11269 & ~w11447;
assign w11449 = ~pi019 & w11246;
assign w11450 = w11442 & ~w11449;
assign w11451 = ~w11448 & w11450;
assign w11452 = ~w11333 & w11451;
assign w11453 = pi023 & w11440;
assign w11454 = pi022 & w11411;
assign w11455 = pi020 & w11387;
assign w11456 = pi021 & w11366;
assign w11457 = ~w11453 & ~w11454;
assign w11458 = ~w11455 & ~w11456;
assign w11459 = w11457 & w11458;
assign w11460 = w10808 & w11459;
assign w11461 = ~w11452 & w11460;
assign w11462 = ~w10809 & ~w11461;
assign w11463 = w10549 & ~w10629;
assign w11464 = (w10929 & ~w11265) | (w10929 & w16712) | (~w11265 & w16712);
assign w11465 = (w10812 & ~w11322) | (w10812 & w18421) | (~w11322 & w18421);
assign w11466 = (w11000 & ~w11157) | (w11000 & w18422) | (~w11157 & w18422);
assign w11467 = (w10552 & ~w11101) | (w10552 & w17320) | (~w11101 & w17320);
assign w11468 = w8499 & ~w11048;
assign w11469 = w6464 & ~w10811;
assign w11470 = w5431 & ~w10903;
assign w11471 = ~w11469 & ~w11470;
assign w11472 = ~w11468 & w11471;
assign w11473 = ~w11467 & w11472;
assign w11474 = ~w11466 & w11473;
assign w11475 = ~w11465 & w11474;
assign w11476 = ~w11464 & w11475;
assign w11477 = (w10550 & ~w11410) | (w10550 & w16713) | (~w11410 & w16713);
assign w11478 = (w10551 & ~w11386) | (w10551 & w16714) | (~w11386 & w16714);
assign w11479 = ~w11477 & ~w11478;
assign w11480 = w11476 & w11479;
assign w11481 = ~w11463 & w11480;
assign w11482 = (~w10532 & ~w10568) | (~w10532 & w18423) | (~w10568 & w18423);
assign w11483 = w11481 & ~w11482;
assign w11484 = ~w5158 & w18483;
assign w11485 = w10574 & ~w10899;
assign w11486 = ~w10899 & w17321;
assign w11487 = (w10580 & ~w11142) | (w10580 & w16716) | (~w11142 & w16716);
assign w11488 = ~w6036 & w11487;
assign w11489 = w10514 & ~w11306;
assign w11490 = ~w11306 & w17322;
assign w11491 = (w10545 & ~w10987) | (w10545 & w16717) | (~w10987 & w16717);
assign w11492 = (~w10987 & w17323) | (~w10987 & w17324) | (w17323 & w17324);
assign w11493 = w9015 & w10944;
assign w11494 = w10924 & w11493;
assign w11495 = (w10572 & ~w10924) | (w10572 & w16718) | (~w10924 & w16718);
assign w11496 = (~w10924 & w17325) | (~w10924 & w17326) | (w17325 & w17326);
assign w11497 = (w10578 & ~w10852) | (w10578 & w16719) | (~w10852 & w16719);
assign w11498 = (~w10852 & w17327) | (~w10852 & w17328) | (w17327 & w17328);
assign w11499 = (~w10542 & ~w10604) | (~w10542 & w17329) | (~w10604 & w17329);
assign w11500 = ~w10386 & w11499;
assign w11501 = (w10576 & ~w11041) | (w10576 & w16720) | (~w11041 & w16720);
assign w11502 = ~w3860 & w11501;
assign w11503 = (w10586 & ~w11089) | (w10586 & w16721) | (~w11089 & w16721);
assign w11504 = ~w4687 & w11503;
assign w11505 = w6467 & w8479;
assign w11506 = ~w8548 & w11505;
assign w11507 = ~w4280 & w11506;
assign w11508 = w11503 & w18424;
assign w11509 = (w10512 & ~w11244) | (w10512 & w16722) | (~w11244 & w16722);
assign w11510 = w10672 & ~w10705;
assign w11511 = ~w10804 & ~w11510;
assign w11512 = (w10520 & ~w11364) | (w10520 & w16723) | (~w11364 & w16723);
assign w11513 = ~w8172 & w11512;
assign w11514 = ~w9672 & ~w11440;
assign w11515 = ~w11440 & w17330;
assign w11516 = w10772 & w11511;
assign w11517 = (w11516 & ~w11509) | (w11516 & w17331) | (~w11509 & w17331);
assign w11518 = ~w11513 & ~w11515;
assign w11519 = w11517 & w11518;
assign w11520 = ~w11484 & ~w11486;
assign w11521 = ~w11488 & ~w11490;
assign w11522 = ~w11492 & ~w11496;
assign w11523 = ~w11498 & ~w11500;
assign w11524 = ~w11502 & w11523;
assign w11525 = w11521 & w11522;
assign w11526 = w11519 & w17332;
assign w11527 = w11524 & w11525;
assign w11528 = w11526 & w11527;
assign w11529 = w11483 & w11528;
assign w11530 = ~w532 & w11495;
assign w11531 = ~w5918 & w11487;
assign w11532 = ~w1546 & w11491;
assign w11533 = ~w5071 & w18483;
assign w11534 = ~w10415 & w11499;
assign w11535 = ~w3773 & w11501;
assign w11536 = ~w1917 & w11485;
assign w11537 = ~w4192 & w9345;
assign w11538 = w11503 & w11537;
assign w11539 = ~w6724 & w11489;
assign w11540 = (w16722 & w18425) | (w16722 & w18426) | (w18425 & w18426);
assign w11541 = ~w3139 & w11497;
assign w11542 = ~w8777 & ~w9005;
assign w11543 = ~w11440 & w17333;
assign w11544 = (~w11511 & ~w11512) | (~w11511 & w17334) | (~w11512 & w17334);
assign w11545 = ~w11540 & ~w11543;
assign w11546 = w11544 & w11545;
assign w11547 = ~w11530 & ~w11531;
assign w11548 = ~w11532 & ~w11533;
assign w11549 = ~w11534 & ~w11535;
assign w11550 = ~w11536 & ~w11538;
assign w11551 = ~w11539 & ~w11541;
assign w11552 = w11550 & w11551;
assign w11553 = w11548 & w11549;
assign w11554 = w11546 & w11547;
assign w11555 = w11553 & w11554;
assign w11556 = w11552 & w11555;
assign w11557 = (pi027 & ~w11555) | (pi027 & w17335) | (~w11555 & w17335);
assign w11558 = w11529 & w11557;
assign w11559 = w11483 & w11556;
assign w11560 = pi028 & w11559;
assign w11561 = ~w950 & w4729;
assign w11562 = ~w10671 & w11561;
assign w11563 = w2627 & w11562;
assign w11564 = w6099 & w11563;
assign w11565 = w10335 & w11564;
assign w11566 = w10313 & w11565;
assign w11567 = w10682 & w11566;
assign w11568 = pi264 & ~pi272;
assign w11569 = pi263 & ~pi271;
assign w11570 = ~pi264 & pi272;
assign w11571 = ~pi265 & pi273;
assign w11572 = pi265 & ~pi273;
assign w11573 = pi266 & ~pi274;
assign w11574 = ~pi266 & pi274;
assign w11575 = ~pi267 & pi275;
assign w11576 = pi269 & ~pi277;
assign w11577 = ~pi269 & pi277;
assign w11578 = pi270 & ~pi278;
assign w11579 = ~w11577 & w11578;
assign w11580 = ~w11576 & ~w11579;
assign w11581 = ~pi276 & ~w11580;
assign w11582 = pi267 & ~pi275;
assign w11583 = pi276 & w11580;
assign w11584 = pi268 & ~w11583;
assign w11585 = ~w11581 & ~w11582;
assign w11586 = ~w11584 & w11585;
assign w11587 = ~w11574 & ~w11575;
assign w11588 = ~w11586 & w11587;
assign w11589 = ~w11572 & ~w11573;
assign w11590 = ~w11588 & w11589;
assign w11591 = ~w11570 & ~w11571;
assign w11592 = ~w11590 & w11591;
assign w11593 = ~w11568 & ~w11569;
assign w11594 = ~w11592 & w11593;
assign w11595 = ~w1671 & ~w6814;
assign w11596 = w9577 & w11595;
assign w11597 = pi247 & pi263;
assign w11598 = w10683 & w11597;
assign w11599 = ~pi271 & ~w957;
assign w11600 = ~w10644 & w11599;
assign w11601 = ~w11598 & ~w11600;
assign w11602 = w10673 & w10691;
assign w11603 = ~pi271 & ~w112;
assign w11604 = w7997 & w11603;
assign w11605 = ~w10674 & w11604;
assign w11606 = ~w11602 & ~w11605;
assign w11607 = w9571 & w9619;
assign w11608 = w11596 & w11607;
assign w11609 = ~w11601 & w11608;
assign w11610 = w5398 & w10686;
assign w11611 = ~w11606 & w11610;
assign w11612 = w562 & w11609;
assign w11613 = ~w2101 & w8960;
assign w11614 = w11612 & w11613;
assign w11615 = ~w1451 & w11611;
assign w11616 = w11614 & w11615;
assign w11617 = ~w3252 & ~w4953;
assign w11618 = ~w5888 & ~w6782;
assign w11619 = w9600 & ~w10443;
assign w11620 = w10695 & ~w10741;
assign w11621 = w11619 & w11620;
assign w11622 = w11617 & w11618;
assign w11623 = ~w3886 & w11616;
assign w11624 = w11622 & w11623;
assign w11625 = ~w4249 & w11621;
assign w11626 = w10322 & ~w11594;
assign w11627 = w11625 & w11626;
assign w11628 = ~w7465 & w11624;
assign w11629 = w11627 & w11628;
assign w11630 = w8084 & w8806;
assign w11631 = w10642 & w11630;
assign w11632 = w11629 & w11631;
assign w11633 = w11567 & w11632;
assign w11634 = w10330 & w11633;
assign w11635 = w8999 & w11634;
assign w11636 = pi030 & w11635;
assign w11637 = ~pi255 & ~pi263;
assign w11638 = pi167 & w5346;
assign w11639 = w6108 & w11638;
assign w11640 = pi263 & ~w11639;
assign w11641 = pi247 & w10673;
assign w11642 = ~w11640 & w11641;
assign w11643 = ~w11637 & ~w11642;
assign w11644 = ~pi263 & pi271;
assign w11645 = ~w11594 & ~w11644;
assign w11646 = ~w1849 & w1852;
assign w11647 = w1829 & ~w11646;
assign w11648 = ~w957 & w4730;
assign w11649 = w10319 & w11648;
assign w11650 = w4056 & w11596;
assign w11651 = w11649 & w11650;
assign w11652 = w8002 & w11651;
assign w11653 = w593 & w11652;
assign w11654 = w1482 & w11653;
assign w11655 = w10339 & ~w11643;
assign w11656 = w11654 & w11655;
assign w11657 = ~w2812 & ~w3916;
assign w11658 = ~w6811 & w9600;
assign w11659 = ~w10472 & ~w11647;
assign w11660 = w11658 & w11659;
assign w11661 = w11656 & w11657;
assign w11662 = w4983 & w10697;
assign w11663 = w11661 & w11662;
assign w11664 = ~w4220 & w11660;
assign w11665 = ~w6006 & ~w10770;
assign w11666 = w11664 & w11665;
assign w11667 = w10641 & w11663;
assign w11668 = ~w11645 & w11667;
assign w11669 = w8835 & w11666;
assign w11670 = w11668 & w11669;
assign w11671 = ~w8113 & w11670;
assign w11672 = ~w7436 & w11671;
assign w11673 = w11567 & w11672;
assign w11674 = w10332 & w11673;
assign w11675 = w8999 & w11674;
assign w11676 = pi029 & w11675;
assign w11677 = ~w11636 & ~w11676;
assign w11678 = ~w11558 & w11677;
assign w11679 = ~w11560 & w11678;
assign w11680 = ~w11440 & w18427;
assign w11681 = ~w10478 & w11499;
assign w11682 = (w10521 & ~w11364) | (w10521 & w17336) | (~w11364 & w17336);
assign w11683 = (w10531 & ~w10852) | (w10531 & w17337) | (~w10852 & w17337);
assign w11684 = ~w10052 & ~w10899;
assign w11685 = w10518 & w11684;
assign w11686 = w10515 & ~w11306;
assign w11687 = (w10548 & ~w11142) | (w10548 & w17338) | (~w11142 & w17338);
assign w11688 = (w16722 & w18428) | (w16722 & w18429) | (w18428 & w18429);
assign w11689 = (w10526 & ~w11089) | (w10526 & w18430) | (~w11089 & w18430);
assign w11690 = (w10517 & ~w11041) | (w10517 & w17339) | (~w11041 & w17339);
assign w11691 = (w10546 & ~w10987) | (w10546 & w17340) | (~w10987 & w17340);
assign w11692 = (w10523 & ~w11195) | (w10523 & w17341) | (~w11195 & w17341);
assign w11693 = w10529 & ~w11494;
assign w11694 = w11482 & ~w11682;
assign w11695 = ~w11680 & w11694;
assign w11696 = ~w11683 & ~w11686;
assign w11697 = ~w11687 & ~w11688;
assign w11698 = ~w11689 & ~w11690;
assign w11699 = ~w11691 & ~w11692;
assign w11700 = ~w11693 & w11699;
assign w11701 = w11697 & w11698;
assign w11702 = w11695 & w11696;
assign w11703 = ~w11681 & ~w11685;
assign w11704 = w11702 & w11703;
assign w11705 = w11700 & w11701;
assign w11706 = w11704 & w11705;
assign w11707 = w11481 & w11706;
assign w11708 = ~pi026 & w11707;
assign w11709 = (w10577 & ~w11041) | (w10577 & w17342) | (~w11041 & w17342);
assign w11710 = w10415 & ~w10705;
assign w11711 = w10386 & ~w10804;
assign w11712 = (w10585 & ~w11364) | (w10585 & w17343) | (~w11364 & w17343);
assign w11713 = (w10583 & ~w11244) | (w10583 & w17344) | (~w11244 & w17344);
assign w11714 = w10575 & ~w10899;
assign w11715 = w154 & w11495;
assign w11716 = w10584 & ~w11306;
assign w11717 = (w10582 & ~w10987) | (w10582 & w17345) | (~w10987 & w17345);
assign w11718 = (w10581 & ~w11142) | (w10581 & w17346) | (~w11142 & w17346);
assign w11719 = (w10588 & ~w11089) | (w10588 & w18431) | (~w11089 & w18431);
assign w11720 = (w10579 & ~w10852) | (w10579 & w17347) | (~w10852 & w17347);
assign w11721 = w10478 & w11482;
assign w11722 = (w10571 & ~w11195) | (w10571 & w17348) | (~w11195 & w17348);
assign w11723 = w10474 & ~w11710;
assign w11724 = ~w11711 & w11723;
assign w11725 = (w11724 & w11440) | (w11724 & w18432) | (w11440 & w18432);
assign w11726 = ~w11712 & ~w11713;
assign w11727 = w11725 & w11726;
assign w11728 = w11499 & ~w11709;
assign w11729 = ~w11714 & ~w11716;
assign w11730 = ~w11717 & ~w11718;
assign w11731 = ~w11719 & ~w11720;
assign w11732 = ~w11721 & ~w11722;
assign w11733 = w11731 & w11732;
assign w11734 = w11729 & w11730;
assign w11735 = w11727 & w18433;
assign w11736 = w11733 & w11734;
assign w11737 = w11735 & w11736;
assign w11738 = w11481 & w11737;
assign w11739 = ~w10899 & w17349;
assign w11740 = w10250 & w11503;
assign w11741 = (w10607 & ~w11195) | (w10607 & w16724) | (~w11195 & w16724);
assign w11742 = w10616 & ~w11306;
assign w11743 = w10247 & w11514;
assign w11744 = (~w9730 & ~w11364) | (~w9730 & w16725) | (~w11364 & w16725);
assign w11745 = w10249 & w11744;
assign w11746 = (~w10130 & ~w10924) | (~w10130 & w16726) | (~w10924 & w16726);
assign w11747 = w10258 & w11746;
assign w11748 = (~w10987 & w17350) | (~w10987 & w17351) | (w17350 & w17351);
assign w11749 = ~w5709 & w11487;
assign w11750 = (~w11041 & w17352) | (~w11041 & w17353) | (w17352 & w17353);
assign w11751 = (~w10852 & w17354) | (~w10852 & w17355) | (w17354 & w17355);
assign w11752 = w7288 & w11509;
assign w11753 = w11463 & ~w11741;
assign w11754 = ~w11742 & ~w11743;
assign w11755 = ~w11745 & ~w11752;
assign w11756 = w11754 & w11755;
assign w11757 = ~w11739 & w11753;
assign w11758 = ~w11740 & ~w11747;
assign w11759 = ~w11748 & ~w11749;
assign w11760 = ~w11750 & ~w11751;
assign w11761 = w11759 & w11760;
assign w11762 = w11757 & w11758;
assign w11763 = w11756 & w11762;
assign w11764 = w11480 & w11761;
assign w11765 = w11763 & w11764;
assign w11766 = ~w11738 & ~w11765;
assign w11767 = w11763 & w17356;
assign w11768 = pi025 & w11738;
assign w11769 = ~w11707 & ~w11767;
assign w11770 = ~w11768 & w11769;
assign w11771 = ~w11766 & w11770;
assign w11772 = ~pi027 & w11529;
assign w11773 = ~w11559 & ~w11708;
assign w11774 = ~w11772 & w11773;
assign w11775 = ~w11771 & w11774;
assign w11776 = w11679 & ~w11775;
assign w11777 = (~w10924 & w17357) | (~w10924 & w17358) | (w17357 & w17358);
assign w11778 = ~w10899 & w10973;
assign w11779 = (w10953 & ~w11386) | (w10953 & w16727) | (~w11386 & w16727);
assign w11780 = (w10972 & ~w10628) | (w10972 & w17816) | (~w10628 & w17816);
assign w11781 = (w16722 & w17817) | (w16722 & w17818) | (w17817 & w17818);
assign w11782 = (w16725 & w17819) | (w16725 & w17820) | (w17819 & w17820);
assign w11783 = (w10951 & ~w10852) | (w10951 & w16728) | (~w10852 & w16728);
assign w11784 = (w10970 & ~w11195) | (w10970 & w17359) | (~w11195 & w17359);
assign w11785 = (w10967 & ~w11142) | (w10967 & w17360) | (~w11142 & w17360);
assign w11786 = w1755 & w11477;
assign w11787 = w10950 & ~w11440;
assign w11788 = ~w10605 & w10956;
assign w11789 = ~w11779 & ~w11780;
assign w11790 = ~w11787 & w11789;
assign w11791 = ~w11778 & ~w11781;
assign w11792 = ~w11782 & ~w11783;
assign w11793 = ~w11784 & ~w11785;
assign w11794 = ~w11786 & ~w11788;
assign w11795 = w11793 & w11794;
assign w11796 = w11791 & w11792;
assign w11797 = ~w11777 & w11790;
assign w11798 = w11796 & w11797;
assign w11799 = w11795 & w11798;
assign w11800 = (w10975 & ~w11041) | (w10975 & w16729) | (~w11041 & w16729);
assign w11801 = w10949 & ~w11103;
assign w11802 = (w10954 & ~w11157) | (w10954 & w18434) | (~w11157 & w18434);
assign w11803 = (w4808 & ~w10120) | (w4808 & w17361) | (~w10120 & w17361);
assign w11804 = w6317 & ~w10811;
assign w11805 = w7920 & ~w11048;
assign w11806 = w1546 & ~w10705;
assign w11807 = w1515 & ~w10804;
assign w11808 = w10966 & ~w11323;
assign w11809 = w10965 & ~w11306;
assign w11810 = (w10976 & ~w11089) | (w10976 & w16730) | (~w11089 & w16730);
assign w11811 = w1137 & w11464;
assign w11812 = ~w10569 & w10955;
assign w11813 = w1484 & ~w3346;
assign w11814 = ~w11806 & w11813;
assign w11815 = ~w11807 & w11814;
assign w11816 = ~w11803 & w11815;
assign w11817 = ~w11805 & w11816;
assign w11818 = ~w11804 & w11817;
assign w11819 = ~w11802 & w11818;
assign w11820 = ~w11801 & w11819;
assign w11821 = ~w11808 & w11820;
assign w11822 = w11491 & ~w11800;
assign w11823 = ~w11809 & ~w11810;
assign w11824 = ~w11811 & ~w11812;
assign w11825 = w11823 & w11824;
assign w11826 = w11821 & w11822;
assign w11827 = w11825 & w11826;
assign w11828 = w11826 & w17821;
assign w11829 = w11799 & w11828;
assign w11830 = (w10926 & ~w11157) | (w10926 & w18435) | (~w11157 & w18435);
assign w11831 = w6180 & ~w10811;
assign w11832 = w4847 & ~w10903;
assign w11833 = w532 & ~w10705;
assign w11834 = ~w501 & ~w10804;
assign w11835 = w437 & w3346;
assign w11836 = (w10910 & ~w11364) | (w10910 & w16731) | (~w11364 & w16731);
assign w11837 = (w10925 & ~w11322) | (w10925 & w18436) | (~w11322 & w18436);
assign w11838 = (w10933 & ~w10568) | (w10933 & w18437) | (~w10568 & w18437);
assign w11839 = w852 & w11467;
assign w11840 = (w10932 & ~w11386) | (w10932 & w16732) | (~w11386 & w16732);
assign w11841 = (w10906 & ~w11244) | (w10906 & w16733) | (~w11244 & w16733);
assign w11842 = w10907 & ~w10990;
assign w11843 = ~w10185 & ~w11306;
assign w11844 = w10121 & w11843;
assign w11845 = ~w10605 & w10934;
assign w11846 = (~w9882 & ~w11195) | (~w9882 & w16734) | (~w11195 & w16734);
assign w11847 = w10103 & w11846;
assign w11848 = w10927 & ~w11043;
assign w11849 = w659 & w11464;
assign w11850 = w6562 & ~w11835;
assign w11851 = ~w7872 & w11850;
assign w11852 = ~w11833 & w11851;
assign w11853 = ~w11834 & w11852;
assign w11854 = w10892 & w11853;
assign w11855 = ~w11832 & w11854;
assign w11856 = ~w11831 & w11855;
assign w11857 = ~w11830 & w11856;
assign w11858 = ~w11494 & w11857;
assign w11859 = ~w11836 & ~w11837;
assign w11860 = ~w11838 & ~w11839;
assign w11861 = ~w11840 & ~w11841;
assign w11862 = w11860 & w11861;
assign w11863 = w11858 & w11859;
assign w11864 = ~w11842 & ~w11845;
assign w11865 = ~w11848 & ~w11849;
assign w11866 = w11864 & w11865;
assign w11867 = w11862 & w11863;
assign w11868 = ~w11844 & ~w11847;
assign w11869 = w11867 & w11868;
assign w11870 = w11866 & w11869;
assign w11871 = w10908 & ~w11091;
assign w11872 = (w10913 & ~w11142) | (w10913 & w16735) | (~w11142 & w16735);
assign w11873 = (w10911 & ~w10852) | (w10911 & w16736) | (~w10852 & w16736);
assign w11874 = ~w11440 & w18438;
assign w11875 = w10931 & ~w11411;
assign w11876 = ~w10899 & w10904;
assign w11877 = ~w10629 & w10914;
assign w11878 = ~w11875 & ~w11877;
assign w11879 = ~w11871 & w11878;
assign w11880 = ~w11872 & ~w11873;
assign w11881 = ~w11874 & ~w11876;
assign w11882 = w11880 & w11881;
assign w11883 = w11879 & w11882;
assign w11884 = w10947 & w11883;
assign w11885 = w11870 & w11884;
assign w11886 = (w10856 & ~w11089) | (w10856 & w16737) | (~w11089 & w16737);
assign w11887 = (w10893 & ~w10924) | (w10893 & w16738) | (~w10924 & w16738);
assign w11888 = (w10861 & ~w11101) | (w10861 & w17362) | (~w11101 & w17362);
assign w11889 = w6244 & ~w10811;
assign w11890 = w1917 & ~w10705;
assign w11891 = w2260 & w11468;
assign w11892 = (w4797 & ~w10120) | (w4797 & w17363) | (~w10120 & w17363);
assign w11893 = w1886 & ~w10804;
assign w11894 = (w10866 & ~w10852) | (w10866 & w16739) | (~w10852 & w16739);
assign w11895 = (w16725 & w10872) | (w16725 & w17822) | (w10872 & w17822);
assign w11896 = w10013 & w11843;
assign w11897 = w2502 & w11501;
assign w11898 = ~w1825 & w11499;
assign w11899 = (w10891 & ~w11322) | (w10891 & w17364) | (~w11322 & w17364);
assign w11900 = (w10873 & ~w11265) | (w10873 & w16740) | (~w11265 & w16740);
assign w11901 = (w10857 & ~w11386) | (w10857 & w16741) | (~w11386 & w16741);
assign w11902 = (w17365 & ~w10628) | (w17365 & w18439) | (~w10628 & w18439);
assign w11903 = (w10865 & ~w11195) | (w10865 & w17366) | (~w11195 & w17366);
assign w11904 = ~w11440 & w10894;
assign w11905 = (w10869 & ~w11142) | (w10869 & w17367) | (~w11142 & w17367);
assign w11906 = (w10860 & ~w10568) | (w10860 & w17823) | (~w10568 & w17823);
assign w11907 = (w10868 & ~w10987) | (w10868 & w17368) | (~w10987 & w17368);
assign w11908 = (w10870 & ~w11244) | (w10870 & w17369) | (~w11244 & w17369);
assign w11909 = (w10871 & ~w11410) | (w10871 & w17370) | (~w11410 & w17370);
assign w11910 = w2291 & w11466;
assign w11911 = ~w11890 & ~w11893;
assign w11912 = w10049 & w11911;
assign w11913 = (~w10030 & w17371) | (~w10030 & w17372) | (w17371 & w17372);
assign w11914 = ~w11892 & w11913;
assign w11915 = ~w11889 & w11914;
assign w11916 = ~w11891 & w11915;
assign w11917 = ~w11888 & w11916;
assign w11918 = ~w10899 & w11917;
assign w11919 = ~w11899 & ~w11900;
assign w11920 = ~w11901 & ~w11906;
assign w11921 = ~w11908 & w18440;
assign w11922 = w11919 & w11920;
assign w11923 = ~w11886 & w11918;
assign w11924 = ~w11887 & ~w11894;
assign w11925 = ~w11895 & ~w11902;
assign w11926 = ~w11903 & ~w11904;
assign w11927 = ~w11905 & ~w11907;
assign w11928 = w11926 & w11927;
assign w11929 = w11924 & w11925;
assign w11930 = w11922 & w11923;
assign w11931 = ~w11896 & w11921;
assign w11932 = ~w11897 & ~w11898;
assign w11933 = w11931 & w11932;
assign w11934 = w11929 & w11930;
assign w11935 = w11928 & w11934;
assign w11936 = w11933 & w11935;
assign w11937 = (~w11936 & w11885) | (~w11936 & w16742) | (w11885 & w16742);
assign w11938 = w11935 & w17373;
assign w11939 = w4098 & ~w10130;
assign w11940 = ~w11494 & w11939;
assign w11941 = w4092 & w11684;
assign w11942 = w4095 & ~w10990;
assign w11943 = w4096 & ~w11939;
assign w11944 = w4097 & ~w11943;
assign w11945 = ~w11940 & w11944;
assign w11946 = ~w11942 & w11945;
assign w11947 = ~w11941 & w11946;
assign w11948 = ~w11938 & ~w11947;
assign w11949 = ~w11937 & w11948;
assign w11950 = (w11031 & ~w11089) | (w11031 & w16743) | (~w11089 & w16743);
assign w11951 = (w11023 & ~w10987) | (w11023 & w16744) | (~w10987 & w16744);
assign w11952 = (w11009 & ~w11142) | (w11009 & w16745) | (~w11142 & w16745);
assign w11953 = (w11029 & ~w10852) | (w11029 & w16746) | (~w10852 & w16746);
assign w11954 = (w11028 & ~w11244) | (w11028 & w16747) | (~w11244 & w16747);
assign w11955 = w11005 & ~w11102;
assign w11956 = w4038 & w11468;
assign w11957 = w3773 & ~w10705;
assign w11958 = w3860 & ~w10804;
assign w11959 = w11001 & ~w11159;
assign w11960 = (w11003 & ~w10568) | (w11003 & w17824) | (~w10568 & w17824);
assign w11961 = (w11004 & ~w11386) | (w11004 & w16748) | (~w11386 & w16748);
assign w11962 = (w11006 & ~w11322) | (w11006 & w17374) | (~w11322 & w17374);
assign w11963 = w11027 & ~w11440;
assign w11964 = ~w11306 & w11025;
assign w11965 = (w11024 & ~w11364) | (w11024 & w16749) | (~w11364 & w16749);
assign w11966 = ~w10899 & w17375;
assign w11967 = w3830 & w11499;
assign w11968 = (w11008 & ~w11265) | (w11008 & w16750) | (~w11265 & w16750);
assign w11969 = w3449 & w11463;
assign w11970 = (w11007 & ~w11410) | (w11007 & w17376) | (~w11410 & w17376);
assign w11971 = (~w10924 & w17377) | (~w10924 & w17378) | (w17377 & w17378);
assign w11972 = w9957 & w11846;
assign w11973 = w3918 & ~w11957;
assign w11974 = ~w11958 & w11973;
assign w11975 = w10576 & w11974;
assign w11976 = ~w11956 & w11975;
assign w11977 = w11471 & w11976;
assign w11978 = ~w11955 & w11977;
assign w11979 = ~w11959 & w11978;
assign w11980 = ~w11043 & ~w11954;
assign w11981 = ~w11960 & ~w11961;
assign w11982 = ~w11962 & ~w11963;
assign w11983 = ~w11965 & ~w11968;
assign w11984 = ~w11970 & w11983;
assign w11985 = w11981 & w11982;
assign w11986 = w11979 & w11980;
assign w11987 = ~w11950 & ~w11951;
assign w11988 = ~w11952 & ~w11953;
assign w11989 = ~w11969 & w11988;
assign w11990 = w11986 & w11987;
assign w11991 = ~w11964 & ~w11966;
assign w11992 = ~w11967 & ~w11971;
assign w11993 = ~w11972 & w11992;
assign w11994 = w11985 & w18120;
assign w11995 = w11989 & w11990;
assign w11996 = w11995 & w16751;
assign w11997 = (~w10924 & w17379) | (~w10924 & w17380) | (w17379 & w17380);
assign w11998 = w7788 & ~w10899;
assign w11999 = (w7786 & ~w10987) | (w7786 & w16753) | (~w10987 & w16753);
assign w12000 = (w7787 & ~w10852) | (w7787 & w17381) | (~w10852 & w17381);
assign w12001 = w11468 & w11471;
assign w12002 = (w11041 & w17382) | (w11041 & w17383) | (w17382 & w17383);
assign w12003 = ~w11998 & ~w11999;
assign w12004 = ~w12000 & w12003;
assign w12005 = ~w11997 & w12002;
assign w12006 = w12004 & w12005;
assign w12007 = w12004 & w17384;
assign w12008 = (~w10987 & w17385) | (~w10987 & w17386) | (w17385 & w17386);
assign w12009 = (~w10924 & w17387) | (~w10924 & w17388) | (w17387 & w17388);
assign w12010 = (w6266 & ~w10852) | (w6266 & w17389) | (~w10852 & w17389);
assign w12011 = w11469 & ~w11470;
assign w12012 = (w12011 & w10899) | (w12011 & w17390) | (w10899 & w17390);
assign w12013 = ~w12010 & w12012;
assign w12014 = ~w12008 & ~w12009;
assign w12015 = w12013 & w12014;
assign w12016 = ~pi008 & w12015;
assign w12017 = ~w12007 & ~w12016;
assign w12018 = ~w11996 & ~w12017;
assign w12019 = (pi009 & ~w17384) | (pi009 & w18121) | (~w17384 & w18121);
assign w12020 = w11996 & ~w12019;
assign w12021 = ~w12018 & ~w12020;
assign w12022 = w10819 & ~w11306;
assign w12023 = (w10837 & ~w11089) | (w10837 & w16754) | (~w11089 & w16754);
assign w12024 = (w10820 & ~w10924) | (w10820 & w16755) | (~w10924 & w16755);
assign w12025 = (w16725 & w10818) | (w16725 & w18122) | (w10818 & w18122);
assign w12026 = w2873 & w11487;
assign w12027 = ~w11440 & w10829;
assign w12028 = (w10828 & ~w10987) | (w10828 & w16756) | (~w10987 & w16756);
assign w12029 = (w10835 & ~w11195) | (w10835 & w16757) | (~w11195 & w16757);
assign w12030 = (w10817 & ~w11244) | (w10817 & w17391) | (~w11244 & w17391);
assign w12031 = w2931 & w11477;
assign w12032 = ~w11159 & w18123;
assign w12033 = (w10832 & ~w10568) | (w10832 & w18124) | (~w10568 & w18124);
assign w12034 = ~w3019 & w11478;
assign w12035 = w10815 & ~w10899;
assign w12036 = (w10838 & ~w10628) | (w10838 & w18125) | (~w10628 & w18125);
assign w12037 = (w10813 & ~w11322) | (w10813 & w18126) | (~w11322 & w18126);
assign w12038 = (w10836 & ~w11041) | (w10836 & w17392) | (~w11041 & w17392);
assign w12039 = ~w10605 & w10831;
assign w12040 = w10833 & ~w11266;
assign w12041 = (w10830 & ~w11101) | (w10830 & w18127) | (~w11101 & w18127);
assign w12042 = w7797 & ~w10811;
assign w12043 = w7796 & ~w11048;
assign w12044 = w2842 & ~w10803;
assign w12045 = w3139 & ~w10705;
assign w12046 = ~w2813 & ~w3254;
assign w12047 = ~w12044 & w12046;
assign w12048 = ~w12045 & w12047;
assign w12049 = ~w11470 & w12048;
assign w12050 = ~w12043 & w12049;
assign w12051 = ~w12042 & w12050;
assign w12052 = ~w12041 & w12051;
assign w12053 = ~w12030 & w12052;
assign w12054 = ~w12032 & ~w12033;
assign w12055 = ~w12036 & ~w12037;
assign w12056 = ~w12040 & w12055;
assign w12057 = w12053 & w12054;
assign w12058 = w11497 & ~w12022;
assign w12059 = ~w12023 & ~w12024;
assign w12060 = ~w12025 & ~w12027;
assign w12061 = ~w12028 & ~w12029;
assign w12062 = ~w12031 & ~w12034;
assign w12063 = ~w12035 & ~w12038;
assign w12064 = ~w12039 & w12063;
assign w12065 = w12061 & w12062;
assign w12066 = w12059 & w12060;
assign w12067 = w12057 & w12058;
assign w12068 = ~w12026 & w12056;
assign w12069 = w12067 & w12068;
assign w12070 = w12065 & w12066;
assign w12071 = w12064 & w12070;
assign w12072 = w12069 & w12071;
assign w12073 = ~pi006 & w11947;
assign w12074 = ~w12072 & ~w12073;
assign w12075 = w12021 & w12074;
assign w12076 = ~w11949 & w12075;
assign w12077 = w12071 & w17393;
assign w12078 = (~w12015 & ~w16751) | (~w12015 & w17825) | (~w16751 & w17825);
assign w12079 = ~w12077 & w12078;
assign w12080 = w12021 & ~w12079;
assign w12081 = (w16723 & w18128) | (w16723 & w18129) | (w18128 & w18129);
assign w12082 = (w11167 & ~w10924) | (w11167 & w16758) | (~w10924 & w16758);
assign w12083 = ~w10899 & w11172;
assign w12084 = w4895 & w11477;
assign w12085 = (w11176 & ~w11386) | (w11176 & w17394) | (~w11386 & w17394);
assign w12086 = (w11161 & ~w11089) | (w11161 & w16759) | (~w11089 & w16759);
assign w12087 = (w11162 & ~w11244) | (w11162 & w17395) | (~w11244 & w17395);
assign w12088 = ~w12085 & ~w12087;
assign w12089 = ~w12081 & w12088;
assign w12090 = ~w12082 & ~w12083;
assign w12091 = ~w12084 & ~w12086;
assign w12092 = w12090 & w12091;
assign w12093 = w12089 & w12092;
assign w12094 = (w11196 & ~w10852) | (w11196 & w16760) | (~w10852 & w16760);
assign w12095 = (~w10987 & w17396) | (~w10987 & w17397) | (w17396 & w17397);
assign w12096 = (w11169 & ~w11322) | (w11169 & w17398) | (~w11322 & w17398);
assign w12097 = (w11170 & ~w10568) | (w11170 & w17826) | (~w10568 & w17826);
assign w12098 = (w11197 & ~w11142) | (w11197 & w16761) | (~w11142 & w16761);
assign w12099 = (w11173 & ~w11265) | (w11173 & w16762) | (~w11265 & w16762);
assign w12100 = w8466 & w11501;
assign w12101 = w11165 & ~w11306;
assign w12102 = w5071 & ~w10705;
assign w12103 = w5158 & ~w10804;
assign w12104 = (w11164 & ~w10628) | (w11164 & w17827) | (~w10628 & w17827);
assign w12105 = w11198 & ~w11440;
assign w12106 = (w11171 & ~w10604) | (w11171 & w18130) | (~w10604 & w18130);
assign w12107 = ~w12102 & ~w12103;
assign w12108 = w9853 & w12107;
assign w12109 = (w11157 & w18441) | (w11157 & w18442) | (w18441 & w18442);
assign w12110 = w11473 & w12109;
assign w12111 = ~w12096 & ~w12097;
assign w12112 = ~w12099 & ~w12104;
assign w12113 = ~w12105 & w12112;
assign w12114 = w12110 & w12111;
assign w12115 = w11846 & ~w12094;
assign w12116 = ~w12098 & ~w12101;
assign w12117 = ~w12106 & w12116;
assign w12118 = w12114 & w12115;
assign w12119 = ~w12095 & w12113;
assign w12120 = ~w12100 & w12119;
assign w12121 = w12117 & w12118;
assign w12122 = w12120 & w12121;
assign w12123 = w12092 & w17400;
assign w12124 = w12122 & w12123;
assign w12125 = ~w11091 & w11095;
assign w12126 = ~w10899 & w11096;
assign w12127 = w9314 & ~w10990;
assign w12128 = ~w11043 & w11098;
assign w12129 = w9315 & ~w10854;
assign w12130 = w11097 & ~w11494;
assign w12131 = w11467 & w11472;
assign w12132 = ~w12125 & w12131;
assign w12133 = ~w12126 & ~w12127;
assign w12134 = ~w12128 & ~w12129;
assign w12135 = ~w12130 & w12134;
assign w12136 = w12132 & w12133;
assign w12137 = w12135 & w12136;
assign w12138 = ~w12124 & ~w12137;
assign w12139 = (~pi012 & ~w12122) | (~pi012 & w17401) | (~w12122 & w17401);
assign w12140 = ~w12138 & ~w12139;
assign w12141 = (w11059 & ~w11410) | (w11059 & w17402) | (~w11410 & w17402);
assign w12142 = w4313 & w11467;
assign w12143 = (w11069 & ~w11386) | (w11069 & w17403) | (~w11386 & w17403);
assign w12144 = (w11054 & ~w11322) | (w11054 & w18131) | (~w11322 & w18131);
assign w12145 = (w16725 & w11071) | (w16725 & w18132) | (w11071 & w18132);
assign w12146 = w11072 & ~w11159;
assign w12147 = (w11053 & ~w11244) | (w11053 & w17404) | (~w11244 & w17404);
assign w12148 = (w11079 & ~w10628) | (w11079 & w18133) | (~w10628 & w18133);
assign w12149 = (w11073 & ~w10852) | (w11073 & w16763) | (~w10852 & w16763);
assign w12150 = (w11078 & ~w11195) | (w11078 & w16764) | (~w11195 & w16764);
assign w12151 = (w11052 & ~w11041) | (w11052 & w16765) | (~w11041 & w16765);
assign w12152 = ~w1292 & w11491;
assign w12153 = (w11075 & ~w11142) | (w11075 & w16766) | (~w11142 & w16766);
assign w12154 = (w11074 & ~w10924) | (w11074 & w16767) | (~w10924 & w16767);
assign w12155 = w11077 & ~w11306;
assign w12156 = ~w4400 & w11464;
assign w12157 = w4280 & ~w10804;
assign w12158 = w4192 & ~w10705;
assign w12159 = ~w10899 & w11070;
assign w12160 = w9904 & w11514;
assign w12161 = ~w10605 & w11058;
assign w12162 = ~w10569 & w11056;
assign w12163 = w4251 & ~w12158;
assign w12164 = ~w12157 & w12163;
assign w12165 = w11506 & w12164;
assign w12166 = w11472 & w12165;
assign w12167 = ~w12146 & w12166;
assign w12168 = ~w12141 & ~w12142;
assign w12169 = ~w12143 & ~w12144;
assign w12170 = ~w12147 & ~w12148;
assign w12171 = ~w12162 & w12170;
assign w12172 = w12168 & w12169;
assign w12173 = ~w12145 & w12167;
assign w12174 = ~w12149 & ~w12150;
assign w12175 = ~w12151 & ~w12153;
assign w12176 = ~w12154 & ~w12155;
assign w12177 = ~w12156 & ~w12159;
assign w12178 = ~w12160 & ~w12161;
assign w12179 = w12177 & w12178;
assign w12180 = w12175 & w12176;
assign w12181 = w12173 & w12174;
assign w12182 = w12171 & w12172;
assign w12183 = w11504 & ~w12152;
assign w12184 = w12182 & w12183;
assign w12185 = w12180 & w12181;
assign w12186 = w12179 & w12185;
assign w12187 = w12184 & w12186;
assign w12188 = pi010 & w12006;
assign w12189 = ~w12187 & ~w12188;
assign w12190 = ~w12140 & w12189;
assign w12191 = ~w12080 & w12190;
assign w12192 = ~w12076 & w12191;
assign w12193 = (~w12137 & ~w17405) | (~w12137 & w18134) | (~w17405 & w18134);
assign w12194 = ~w12140 & ~w12193;
assign w12195 = (w11121 & ~w10604) | (w11121 & w17406) | (~w10604 & w17406);
assign w12196 = (w11106 & ~w11410) | (w11106 & w16768) | (~w11410 & w16768);
assign w12197 = w11105 & ~w11306;
assign w12198 = (w11129 & ~w11089) | (w11129 & w16769) | (~w11089 & w16769);
assign w12199 = (w11110 & ~w11041) | (w11110 & w16770) | (~w11041 & w16770);
assign w12200 = (w11109 & ~w10852) | (w11109 & w17407) | (~w10852 & w17407);
assign w12201 = w11124 & ~w11440;
assign w12202 = ~w10569 & w11120;
assign w12203 = ~w12196 & ~w12201;
assign w12204 = ~w12202 & w12203;
assign w12205 = ~w12195 & ~w12197;
assign w12206 = ~w12198 & ~w12199;
assign w12207 = ~w12200 & w12206;
assign w12208 = w12204 & w12205;
assign w12209 = w12207 & w12208;
assign w12210 = ~w10899 & w11126;
assign w12211 = ~w1329 & w11491;
assign w12212 = w6098 & w11465;
assign w12213 = (w11119 & ~w11195) | (w11119 & w17408) | (~w11195 & w17408);
assign w12214 = (w11111 & ~w10924) | (w11111 & w17409) | (~w10924 & w17409);
assign w12215 = w5709 & w11463;
assign w12216 = w5918 & ~w10705;
assign w12217 = w6036 & ~w10804;
assign w12218 = (w11125 & ~w11244) | (w11125 & w16772) | (~w11244 & w16772);
assign w12219 = (w11128 & ~w11386) | (w11128 & w16773) | (~w11386 & w16773);
assign w12220 = (w11107 & ~w11364) | (w11107 & w17410) | (~w11364 & w17410);
assign w12221 = ~w6007 & ~w12216;
assign w12222 = ~w12217 & w12221;
assign w12223 = (w11265 & w17411) | (w11265 & w17412) | (w17411 & w17412);
assign w12224 = ~w12218 & ~w12219;
assign w12225 = ~w12220 & w12224;
assign w12226 = w11474 & w12223;
assign w12227 = w11487 & ~w12210;
assign w12228 = ~w12212 & ~w12213;
assign w12229 = ~w12214 & ~w12215;
assign w12230 = w12228 & w12229;
assign w12231 = w12226 & w12227;
assign w12232 = ~w12211 & w12225;
assign w12233 = w12231 & w12232;
assign w12234 = w12230 & w12233;
assign w12235 = w12208 & w17828;
assign w12236 = w12234 & w12235;
assign w12237 = ~w10899 & w17413;
assign w12238 = (~w10987 & w17414) | (~w10987 & w17415) | (w17414 & w17415);
assign w12239 = w9832 & w11846;
assign w12240 = (w11151 & ~w11089) | (w11151 & w16774) | (~w11089 & w16774);
assign w12241 = (w11150 & ~w10852) | (w11150 & w17416) | (~w10852 & w17416);
assign w12242 = (w11148 & ~w11041) | (w11148 & w17417) | (~w11041 & w17417);
assign w12243 = w11145 & ~w11494;
assign w12244 = w11466 & w11473;
assign w12245 = ~w12240 & w12244;
assign w12246 = ~w12241 & ~w12242;
assign w12247 = ~w12243 & w12246;
assign w12248 = ~w12237 & w12245;
assign w12249 = ~w12238 & ~w12239;
assign w12250 = w12248 & w12249;
assign w12251 = w12247 & w12250;
assign w12252 = (~w12251 & ~w12234) | (~w12251 & w17829) | (~w12234 & w17829);
assign w12253 = w9164 & w11503;
assign w12254 = ~w10899 & w11309;
assign w12255 = (w11310 & ~w10987) | (w11310 & w16775) | (~w10987 & w16775);
assign w12256 = (w11313 & ~w11142) | (w11313 & w16776) | (~w11142 & w16776);
assign w12257 = (~w10924 & w17418) | (~w10924 & w17419) | (w17418 & w17419);
assign w12258 = ~w5224 & w18483;
assign w12259 = (w11311 & ~w10852) | (w11311 & w16777) | (~w10852 & w16777);
assign w12260 = ~w3683 & w11501;
assign w12261 = w11465 & w11474;
assign w12262 = ~w12254 & ~w12255;
assign w12263 = ~w12256 & ~w12259;
assign w12264 = w12262 & w12263;
assign w12265 = ~w12253 & w12261;
assign w12266 = ~w12257 & ~w12258;
assign w12267 = ~w12260 & w12266;
assign w12268 = w12264 & w12265;
assign w12269 = w12267 & w12268;
assign w12270 = w12268 & w17420;
assign w12271 = (w11286 & ~w11195) | (w11286 & w16778) | (~w11195 & w16778);
assign w12272 = w6999 & w11478;
assign w12273 = (~w10924 & w17915) | (~w10924 & w17916) | (w17915 & w17916);
assign w12274 = (w11287 & ~w10987) | (w11287 & w16779) | (~w10987 & w16779);
assign w12275 = w6871 & w11499;
assign w12276 = (w11271 & ~w11142) | (w11271 & w16780) | (~w11142 & w16780);
assign w12277 = ~w10899 & w11274;
assign w12278 = (w11275 & ~w10852) | (w11275 & w16781) | (~w10852 & w16781);
assign w12279 = (w11276 & ~w11089) | (w11276 & w16782) | (~w11089 & w16782);
assign w12280 = (w11285 & ~w10568) | (w11285 & w18135) | (~w10568 & w18135);
assign w12281 = (w11280 & ~w11265) | (w11280 & w16783) | (~w11265 & w16783);
assign w12282 = (w11277 & ~w11410) | (w11277 & w16784) | (~w11410 & w16784);
assign w12283 = (w11281 & ~w11244) | (w11281 & w16785) | (~w11244 & w16785);
assign w12284 = (w11278 & ~w11364) | (w11278 & w16786) | (~w11364 & w16786);
assign w12285 = w7962 & w11501;
assign w12286 = ~w10629 & w11282;
assign w12287 = w6724 & ~w10705;
assign w12288 = w6753 & ~w10804;
assign w12289 = w6813 & ~w12287;
assign w12290 = ~w12288 & w12289;
assign w12291 = (w12290 & w11440) | (w12290 & w17421) | (w11440 & w17421);
assign w12292 = ~w12281 & ~w12282;
assign w12293 = ~w12283 & ~w12284;
assign w12294 = w11489 & w12291;
assign w12295 = ~w12271 & ~w12272;
assign w12296 = ~w12274 & ~w12276;
assign w12297 = ~w12277 & ~w12278;
assign w12298 = ~w12279 & ~w12280;
assign w12299 = ~w12286 & w12298;
assign w12300 = w12296 & w12297;
assign w12301 = w12294 & w12295;
assign w12302 = w12293 & w18443;
assign w12303 = ~w12273 & ~w12275;
assign w12304 = ~w12285 & w12303;
assign w12305 = w12301 & w12302;
assign w12306 = w12299 & w12300;
assign w12307 = w12305 & w17830;
assign w12308 = ~w12270 & ~w12307;
assign w12309 = ~pi013 & w12124;
assign w12310 = ~w1168 & w11491;
assign w12311 = ~w10899 & w11370;
assign w12312 = (w11376 & ~w11244) | (w11376 & w16787) | (~w11244 & w16787);
assign w12313 = w3019 & w11497;
assign w12314 = (w11371 & ~w11195) | (w11371 & w16788) | (~w11195 & w16788);
assign w12315 = (w11369 & ~w11041) | (w11369 & w16789) | (~w11041 & w16789);
assign w12316 = w9741 & w11746;
assign w12317 = (w11374 & ~w11142) | (w11374 & w16790) | (~w11142 & w16790);
assign w12318 = ~w11306 & w11375;
assign w12319 = (w11368 & ~w11089) | (w11368 & w18444) | (~w11089 & w18444);
assign w12320 = w11478 & ~w12312;
assign w12321 = ~w12311 & w12320;
assign w12322 = ~w12314 & ~w12315;
assign w12323 = ~w12317 & ~w12318;
assign w12324 = ~w12319 & w12323;
assign w12325 = w12321 & w12322;
assign w12326 = ~w12310 & ~w12313;
assign w12327 = ~w12316 & w12326;
assign w12328 = w12325 & w17831;
assign w12329 = w12327 & w12328;
assign w12330 = w11475 & w18136;
assign w12331 = ~w10899 & w11341;
assign w12332 = (w11338 & ~w10628) | (w11338 & w17832) | (~w10628 & w17832);
assign w12333 = ~w5738 & w11487;
assign w12334 = w8172 & ~w10804;
assign w12335 = w8143 & ~w10705;
assign w12336 = ~w11306 & w11346;
assign w12337 = (w11339 & ~w11089) | (w11339 & w16791) | (~w11089 & w16791);
assign w12338 = (w11345 & ~w10987) | (w11345 & w16792) | (~w10987 & w16792);
assign w12339 = (w11344 & ~w11195) | (w11344 & w16793) | (~w11195 & w16793);
assign w12340 = (w11340 & ~w10852) | (w11340 & w16794) | (~w10852 & w16794);
assign w12341 = (w11336 & ~w11041) | (w11336 & w16795) | (~w11041 & w16795);
assign w12342 = (w11342 & ~w10604) | (w11342 & w17422) | (~w10604 & w17422);
assign w12343 = (w11343 & ~w10568) | (w11343 & w17833) | (~w10568 & w17833);
assign w12344 = (w11337 & ~w10924) | (w11337 & w16796) | (~w10924 & w16796);
assign w12345 = (w11335 & ~w11410) | (w11335 & w16797) | (~w11410 & w16797);
assign w12346 = w11347 & ~w11440;
assign w12347 = (w16722 & w18137) | (w16722 & w18138) | (w18137 & w18138);
assign w12348 = ~w12334 & ~w12335;
assign w12349 = w9713 & w12348;
assign w12350 = (w16725 & w17834) | (w16725 & w17835) | (w17834 & w17835);
assign w12351 = ~w12332 & ~w12343;
assign w12352 = ~w12345 & ~w12346;
assign w12353 = ~w12331 & w12350;
assign w12354 = ~w12336 & ~w12337;
assign w12355 = ~w12338 & ~w12339;
assign w12356 = ~w12340 & ~w12341;
assign w12357 = ~w12342 & ~w12344;
assign w12358 = ~w12347 & w12357;
assign w12359 = w12355 & w12356;
assign w12360 = w12353 & w12354;
assign w12361 = w12352 & w18445;
assign w12362 = w12360 & w12361;
assign w12363 = w12358 & w12359;
assign w12364 = w12362 & w17836;
assign w12365 = ~w12329 & ~w12364;
assign w12366 = (w17423 & ~w10628) | (w17423 & w18139) | (~w10628 & w18139);
assign w12367 = (w16722 & w17837) | (w16722 & w17838) | (w17837 & w17838);
assign w12368 = w8836 & ~w9005;
assign w12369 = ~w8953 & ~w10804;
assign w12370 = w8777 & ~w10705;
assign w12371 = (w11417 & ~w11041) | (w11417 & w16798) | (~w11041 & w16798);
assign w12372 = (w11415 & ~w11089) | (w11415 & w16799) | (~w11089 & w16799);
assign w12373 = (w11414 & ~w10987) | (w11414 & w16800) | (~w10987 & w16800);
assign w12374 = (w11423 & ~w10568) | (w11423 & w18140) | (~w10568 & w18140);
assign w12375 = (w11412 & ~w11142) | (w11412 & w16801) | (~w11142 & w16801);
assign w12376 = ~w11306 & w11425;
assign w12377 = (w11422 & ~w10604) | (w11422 & w17424) | (~w10604 & w17424);
assign w12378 = (w16725 & w11421) | (w16725 & w17839) | (w11421 & w17839);
assign w12379 = (w11419 & ~w11195) | (w11419 & w16802) | (~w11195 & w16802);
assign w12380 = (w11418 & ~w10852) | (w11418 & w16803) | (~w10852 & w16803);
assign w12381 = (w11413 & ~w10924) | (w11413 & w16804) | (~w10924 & w16804);
assign w12382 = ~w10899 & w11420;
assign w12383 = w12368 & ~w12370;
assign w12384 = ~w12369 & w12383;
assign w12385 = ~w11440 & w17425;
assign w12386 = ~w12366 & w12385;
assign w12387 = ~w12367 & ~w12371;
assign w12388 = ~w12372 & ~w12373;
assign w12389 = ~w12374 & ~w12375;
assign w12390 = ~w12376 & ~w12377;
assign w12391 = ~w12378 & ~w12379;
assign w12392 = ~w12380 & ~w12381;
assign w12393 = ~w12382 & w12392;
assign w12394 = w12390 & w12391;
assign w12395 = w12388 & w12389;
assign w12396 = w12386 & w12387;
assign w12397 = w12395 & w12396;
assign w12398 = w12393 & w12394;
assign w12399 = w12397 & w12398;
assign w12400 = w11480 & w12399;
assign w12401 = (w16722 & w18141) | (w16722 & w18142) | (w18141 & w18142);
assign w12402 = (w11397 & ~w10987) | (w11397 & w16805) | (~w10987 & w16805);
assign w12403 = (w11395 & ~w11089) | (w11395 & w16806) | (~w11089 & w16806);
assign w12404 = (w11394 & ~w11195) | (w11394 & w16807) | (~w11195 & w16807);
assign w12405 = (w11399 & ~w11142) | (w11399 & w16808) | (~w11142 & w16808);
assign w12406 = (w11396 & ~w10924) | (w11396 & w17426) | (~w10924 & w17426);
assign w12407 = ~w11306 & w11392;
assign w12408 = ~w10899 & w11393;
assign w12409 = ~w3534 & w11501;
assign w12410 = (w11390 & ~w11364) | (w11390 & w16809) | (~w11364 & w16809);
assign w12411 = (w11389 & ~w10852) | (w11389 & w16810) | (~w10852 & w16810);
assign w12412 = w11477 & ~w12410;
assign w12413 = ~w12401 & w12412;
assign w12414 = ~w12402 & ~w12403;
assign w12415 = ~w12404 & ~w12405;
assign w12416 = ~w12406 & ~w12407;
assign w12417 = ~w12408 & ~w12411;
assign w12418 = w12416 & w12417;
assign w12419 = w12414 & w12415;
assign w12420 = ~w12409 & w12413;
assign w12421 = w12419 & w12420;
assign w12422 = w12421 & w17427;
assign w12423 = ~w12400 & ~w12422;
assign w12424 = w12365 & w12423;
assign w12425 = ~w7526 & w11499;
assign w12426 = ~w2042 & w11485;
assign w12427 = w9759 & w11746;
assign w12428 = (w11223 & ~w11089) | (w11223 & w16811) | (~w11089 & w16811);
assign w12429 = w7407 & ~w10705;
assign w12430 = (w11221 & ~w10987) | (w11221 & w16812) | (~w10987 & w16812);
assign w12431 = (w11212 & ~w11386) | (w11212 & w16813) | (~w11386 & w16813);
assign w12432 = ~w7495 & ~w10804;
assign w12433 = (w11218 & ~w10568) | (w11218 & w18143) | (~w10568 & w18143);
assign w12434 = w11216 & ~w11306;
assign w12435 = (w11226 & ~w11142) | (w11226 & w16814) | (~w11142 & w16814);
assign w12436 = ~w10629 & w18144;
assign w12437 = (w11219 & ~w11041) | (w11219 & w16815) | (~w11041 & w16815);
assign w12438 = ~w11440 & w11214;
assign w12439 = (w11220 & ~w10852) | (w11220 & w16816) | (~w10852 & w16816);
assign w12440 = w9767 & w11846;
assign w12441 = (w16725 & w18145) | (w16725 & w18146) | (w18145 & w18146);
assign w12442 = w11213 & ~w11411;
assign w12443 = w7466 & ~w12429;
assign w12444 = ~w12432 & w12443;
assign w12445 = (w16722 & w18147) | (w16722 & w18148) | (w18147 & w18148);
assign w12446 = ~w12431 & ~w12433;
assign w12447 = ~w12442 & w12446;
assign w12448 = ~w12428 & w12445;
assign w12449 = ~w12430 & ~w12434;
assign w12450 = ~w12435 & ~w12436;
assign w12451 = ~w12437 & ~w12438;
assign w12452 = ~w12439 & ~w12441;
assign w12453 = w12451 & w12452;
assign w12454 = w12449 & w12450;
assign w12455 = w12447 & w12448;
assign w12456 = ~w12425 & ~w12426;
assign w12457 = ~w12427 & ~w12440;
assign w12458 = w12456 & w12457;
assign w12459 = w12454 & w12455;
assign w12460 = w11476 & w12453;
assign w12461 = w12459 & w12460;
assign w12462 = w12458 & w12461;
assign w12463 = w12461 & w18149;
assign w12464 = ~w10899 & w11248;
assign w12465 = w10212 & w11846;
assign w12466 = ~w11144 & w11247;
assign w12467 = ~w10990 & w11254;
assign w12468 = w9145 & w11503;
assign w12469 = w10217 & w11843;
assign w12470 = ~w2723 & w11497;
assign w12471 = ~w659 & w11495;
assign w12472 = w11464 & w18484;
assign w12473 = ~w12464 & ~w12466;
assign w12474 = ~w12467 & w12473;
assign w12475 = w11475 & w12472;
assign w12476 = ~w12465 & ~w12468;
assign w12477 = ~w12469 & ~w12470;
assign w12478 = ~w12471 & w12477;
assign w12479 = w12475 & w12476;
assign w12480 = w12474 & w12479;
assign w12481 = w12478 & w12480;
assign w12482 = (~pi018 & ~w12461) | (~pi018 & w18150) | (~w12461 & w18150);
assign w12483 = w12481 & w12482;
assign w12484 = w12424 & w18446;
assign w12485 = w12252 & w12308;
assign w12486 = ~w12309 & w12485;
assign w12487 = ~w12194 & w12486;
assign w12488 = w12484 & w12487;
assign w12489 = ~w12192 & w12488;
assign w12490 = w12234 & w17840;
assign w12491 = w12250 & w18447;
assign w12492 = ~w12269 & ~w12491;
assign w12493 = ~w12490 & w12492;
assign w12494 = w12308 & ~w12493;
assign w12495 = ~w12462 & ~w12481;
assign w12496 = pi017 & w12307;
assign w12497 = w12495 & ~w12496;
assign w12498 = ~w12494 & w12497;
assign w12499 = w12484 & ~w12498;
assign w12500 = w12421 & w18151;
assign w12501 = w12328 & w16819;
assign w12502 = w12399 & w16820;
assign w12503 = w12362 & w18152;
assign w12504 = ~w12500 & ~w12501;
assign w12505 = ~w12502 & ~w12503;
assign w12506 = w12504 & w12505;
assign w12507 = w11770 & w12506;
assign w12508 = w11679 & w12507;
assign w12509 = ~w12499 & w12508;
assign w12510 = ~w12489 & w12509;
assign w12511 = ~w11776 & ~w12510;
assign w12512 = ~pi047 & ~w27;
assign w12513 = pi039 & w819;
assign w12514 = w787 & w12513;
assign w12515 = w851 & w12514;
assign w12516 = w3410 & w12515;
assign w12517 = w470 & w12516;
assign w12518 = ~w29 & ~w12517;
assign w12519 = ~w12512 & ~w12518;
assign w12520 = pi048 & w29;
assign w12521 = pi040 & w919;
assign w12522 = ~w12520 & ~w12521;
assign w12523 = pi049 & w29;
assign w12524 = pi041 & w919;
assign w12525 = ~w12523 & ~w12524;
assign w12526 = pi050 & w29;
assign w12527 = pi042 & w919;
assign w12528 = ~w12526 & ~w12527;
assign w12529 = pi051 & w29;
assign w12530 = pi043 & w919;
assign w12531 = ~w12529 & ~w12530;
assign w12532 = pi052 & w29;
assign w12533 = pi044 & w919;
assign w12534 = ~w12532 & ~w12533;
assign w12535 = pi053 & w29;
assign w12536 = pi045 & w919;
assign w12537 = ~w12535 & ~w12536;
assign w12538 = pi054 & w29;
assign w12539 = pi046 & w919;
assign w12540 = ~w12538 & ~w12539;
assign w12541 = pi039 & pi063;
assign w12542 = ~w950 & w12541;
assign w12543 = w922 & w12542;
assign w12544 = ~w1759 & ~w12543;
assign w12545 = pi055 & ~w12544;
assign w12546 = ~w919 & w12517;
assign w12547 = pi047 & w919;
assign w12548 = ~w12546 & ~w12547;
assign w12549 = ~w12545 & w12548;
assign w12550 = pi056 & w1759;
assign w12551 = pi040 & ~w919;
assign w12552 = w918 & w12551;
assign w12553 = pi064 & w955;
assign w12554 = pi048 & w919;
assign w12555 = ~w12550 & ~w12553;
assign w12556 = ~w12554 & w12555;
assign w12557 = ~w12552 & w12556;
assign w12558 = pi057 & w1759;
assign w12559 = pi041 & ~w919;
assign w12560 = w918 & w12559;
assign w12561 = pi065 & w955;
assign w12562 = pi049 & w919;
assign w12563 = ~w12558 & ~w12561;
assign w12564 = ~w12562 & w12563;
assign w12565 = ~w12560 & w12564;
assign w12566 = pi058 & w1759;
assign w12567 = pi042 & ~w919;
assign w12568 = w918 & w12567;
assign w12569 = pi066 & w955;
assign w12570 = pi050 & w919;
assign w12571 = ~w12566 & ~w12569;
assign w12572 = ~w12570 & w12571;
assign w12573 = ~w12568 & w12572;
assign w12574 = pi059 & w1759;
assign w12575 = pi043 & ~w919;
assign w12576 = w918 & w12575;
assign w12577 = pi067 & w955;
assign w12578 = pi051 & w919;
assign w12579 = ~w12574 & ~w12577;
assign w12580 = ~w12578 & w12579;
assign w12581 = ~w12576 & w12580;
assign w12582 = pi060 & w1759;
assign w12583 = pi044 & ~w919;
assign w12584 = w918 & w12583;
assign w12585 = pi068 & w955;
assign w12586 = pi052 & w919;
assign w12587 = ~w12582 & ~w12585;
assign w12588 = ~w12586 & w12587;
assign w12589 = ~w12584 & w12588;
assign w12590 = pi061 & w1759;
assign w12591 = pi045 & ~w919;
assign w12592 = w918 & w12591;
assign w12593 = pi069 & w955;
assign w12594 = pi053 & w919;
assign w12595 = ~w12590 & ~w12593;
assign w12596 = ~w12594 & w12595;
assign w12597 = ~w12592 & w12596;
assign w12598 = pi062 & w1759;
assign w12599 = pi046 & ~w919;
assign w12600 = w918 & w12599;
assign w12601 = pi070 & w955;
assign w12602 = pi054 & w919;
assign w12603 = ~w12598 & ~w12601;
assign w12604 = ~w12602 & w12603;
assign w12605 = ~w12600 & w12604;
assign w12606 = pi071 & w2540;
assign w12607 = ~w918 & w2567;
assign w12608 = w12516 & w12607;
assign w12609 = ~w2564 & w12608;
assign w12610 = pi079 & w6108;
assign w12611 = w2547 & w12610;
assign w12612 = pi063 & w2575;
assign w12613 = pi055 & w1754;
assign w12614 = w2559 & w12613;
assign w12615 = ~w2555 & w12614;
assign w12616 = w3311 & w12615;
assign w12617 = ~w12609 & ~w12611;
assign w12618 = ~w12616 & w12617;
assign w12619 = ~w12606 & ~w12612;
assign w12620 = w12618 & w12619;
assign w12621 = pi072 & w2540;
assign w12622 = pi080 & w2552;
assign w12623 = pi056 & w2562;
assign w12624 = pi040 & w2570;
assign w12625 = pi064 & w2575;
assign w12626 = ~w12621 & ~w12622;
assign w12627 = ~w12623 & ~w12624;
assign w12628 = ~w12625 & w12627;
assign w12629 = w12626 & w12628;
assign w12630 = pi073 & w2540;
assign w12631 = pi081 & w2552;
assign w12632 = pi057 & w2562;
assign w12633 = pi065 & w2575;
assign w12634 = pi041 & w2570;
assign w12635 = ~w12630 & ~w12631;
assign w12636 = ~w12632 & ~w12633;
assign w12637 = ~w12634 & w12636;
assign w12638 = w12635 & w12637;
assign w12639 = pi074 & w2540;
assign w12640 = pi082 & w2552;
assign w12641 = pi058 & w2562;
assign w12642 = pi042 & w2570;
assign w12643 = pi066 & w2575;
assign w12644 = ~w12639 & ~w12640;
assign w12645 = ~w12641 & ~w12642;
assign w12646 = ~w12643 & w12645;
assign w12647 = w12644 & w12646;
assign w12648 = pi075 & w2540;
assign w12649 = pi083 & w2552;
assign w12650 = pi059 & w2562;
assign w12651 = pi067 & w2575;
assign w12652 = pi043 & w2570;
assign w12653 = ~w12648 & ~w12649;
assign w12654 = ~w12650 & ~w12651;
assign w12655 = ~w12652 & w12654;
assign w12656 = w12653 & w12655;
assign w12657 = pi076 & w2540;
assign w12658 = pi084 & w2552;
assign w12659 = pi060 & w2562;
assign w12660 = pi068 & w2575;
assign w12661 = pi044 & w2570;
assign w12662 = ~w12657 & ~w12658;
assign w12663 = ~w12659 & ~w12660;
assign w12664 = ~w12661 & w12663;
assign w12665 = w12662 & w12664;
assign w12666 = pi077 & w2540;
assign w12667 = pi085 & w2552;
assign w12668 = pi061 & w2562;
assign w12669 = pi045 & w2570;
assign w12670 = pi069 & w2575;
assign w12671 = ~w12666 & ~w12667;
assign w12672 = ~w12668 & ~w12669;
assign w12673 = ~w12670 & w12672;
assign w12674 = w12671 & w12673;
assign w12675 = pi078 & w2540;
assign w12676 = pi086 & w2552;
assign w12677 = pi062 & w2562;
assign w12678 = pi046 & w2570;
assign w12679 = pi070 & w2575;
assign w12680 = ~w12675 & ~w12676;
assign w12681 = ~w12677 & ~w12678;
assign w12682 = ~w12679 & w12681;
assign w12683 = w12680 & w12682;
assign w12684 = pi087 & w3296;
assign w12685 = pi063 & w2635;
assign w12686 = pi095 & w2632;
assign w12687 = w1169 & w12613;
assign w12688 = ~w2561 & w12687;
assign w12689 = w3320 & w12688;
assign w12690 = w3309 & w12689;
assign w12691 = pi079 & w2590;
assign w12692 = pi071 & w1948;
assign w12693 = w2386 & ~w3303;
assign w12694 = w3378 & w12693;
assign w12695 = w3302 & w12694;
assign w12696 = w12692 & w12695;
assign w12697 = w3335 & w12516;
assign w12698 = w3330 & w12697;
assign w12699 = ~w12686 & ~w12690;
assign w12700 = ~w12685 & w12699;
assign w12701 = ~w12698 & w12700;
assign w12702 = ~w12684 & ~w12696;
assign w12703 = w12701 & w12702;
assign w12704 = ~w12691 & w12703;
assign w12705 = pi080 & w2590;
assign w12706 = pi096 & w2632;
assign w12707 = pi064 & w2635;
assign w12708 = pi072 & ~w1949;
assign w12709 = w12695 & w12708;
assign w12710 = pi088 & w3296;
assign w12711 = pi056 & w3324;
assign w12712 = pi040 & w3337;
assign w12713 = ~w12706 & ~w12707;
assign w12714 = ~w12711 & w12713;
assign w12715 = ~w12709 & ~w12710;
assign w12716 = ~w12712 & w12715;
assign w12717 = ~w12705 & w12714;
assign w12718 = w12716 & w12717;
assign w12719 = pi081 & w2590;
assign w12720 = pi097 & w2632;
assign w12721 = pi065 & w2635;
assign w12722 = pi041 & w3337;
assign w12723 = pi089 & w3296;
assign w12724 = pi057 & w3324;
assign w12725 = pi073 & ~w1949;
assign w12726 = w12695 & w12725;
assign w12727 = ~w12720 & ~w12721;
assign w12728 = ~w12724 & w12727;
assign w12729 = ~w12722 & ~w12723;
assign w12730 = ~w12726 & w12729;
assign w12731 = ~w12719 & w12728;
assign w12732 = w12730 & w12731;
assign w12733 = pi082 & w2590;
assign w12734 = pi098 & w2632;
assign w12735 = pi066 & w2635;
assign w12736 = pi074 & ~w1949;
assign w12737 = w12695 & w12736;
assign w12738 = pi090 & w3296;
assign w12739 = pi058 & w3324;
assign w12740 = pi042 & w3337;
assign w12741 = ~w12734 & ~w12735;
assign w12742 = ~w12739 & w12741;
assign w12743 = ~w12737 & ~w12738;
assign w12744 = ~w12740 & w12743;
assign w12745 = ~w12733 & w12742;
assign w12746 = w12744 & w12745;
assign w12747 = pi083 & w2590;
assign w12748 = pi099 & w2632;
assign w12749 = pi067 & w2635;
assign w12750 = pi091 & w3296;
assign w12751 = pi043 & w3337;
assign w12752 = pi059 & w3324;
assign w12753 = pi075 & ~w1949;
assign w12754 = w12695 & w12753;
assign w12755 = ~w12748 & ~w12749;
assign w12756 = ~w12752 & w12755;
assign w12757 = ~w12750 & ~w12751;
assign w12758 = ~w12754 & w12757;
assign w12759 = ~w12747 & w12756;
assign w12760 = w12758 & w12759;
assign w12761 = pi084 & w2590;
assign w12762 = pi100 & w2632;
assign w12763 = pi068 & w2635;
assign w12764 = pi076 & ~w1949;
assign w12765 = w12695 & w12764;
assign w12766 = pi092 & w3296;
assign w12767 = pi060 & w3324;
assign w12768 = pi044 & w3337;
assign w12769 = ~w12762 & ~w12763;
assign w12770 = ~w12767 & w12769;
assign w12771 = ~w12765 & ~w12766;
assign w12772 = ~w12768 & w12771;
assign w12773 = ~w12761 & w12770;
assign w12774 = w12772 & w12773;
assign w12775 = pi085 & w2590;
assign w12776 = pi101 & w2632;
assign w12777 = pi069 & w2635;
assign w12778 = pi045 & w3337;
assign w12779 = pi077 & ~w1949;
assign w12780 = w12695 & w12779;
assign w12781 = pi061 & w3324;
assign w12782 = pi093 & w3296;
assign w12783 = ~w12776 & ~w12777;
assign w12784 = ~w12781 & w12783;
assign w12785 = ~w12778 & ~w12780;
assign w12786 = ~w12782 & w12785;
assign w12787 = ~w12775 & w12784;
assign w12788 = w12786 & w12787;
assign w12789 = pi086 & w2590;
assign w12790 = pi102 & w2632;
assign w12791 = pi070 & w2635;
assign w12792 = pi078 & ~w1949;
assign w12793 = w12695 & w12792;
assign w12794 = pi094 & w3296;
assign w12795 = pi062 & w3324;
assign w12796 = pi046 & w3337;
assign w12797 = ~w12790 & ~w12791;
assign w12798 = ~w12795 & w12797;
assign w12799 = ~w12793 & ~w12794;
assign w12800 = ~w12796 & w12799;
assign w12801 = ~w12789 & w12798;
assign w12802 = w12800 & w12801;
assign w12803 = pi039 & pi111;
assign w12804 = w4069 & w12803;
assign w12805 = pi095 & w4083;
assign w12806 = pi079 & w3353;
assign w12807 = pi103 & w4051;
assign w12808 = pi087 & w3137;
assign w12809 = w3165 & w12808;
assign w12810 = w3111 & w12809;
assign w12811 = w3256 & w12810;
assign w12812 = w3285 & w12811;
assign w12813 = ~w3389 & w12812;
assign w12814 = w3399 & w12813;
assign w12815 = pi039 & pi127;
assign w12816 = ~w849 & w12815;
assign w12817 = w5594 & w12816;
assign w12818 = w3419 & w12817;
assign w12819 = pi055 & w4094;
assign w12820 = w3375 & w3385;
assign w12821 = w12692 & w12820;
assign w12822 = ~w12804 & ~w12807;
assign w12823 = ~w12814 & ~w12818;
assign w12824 = w12822 & w12823;
assign w12825 = ~w12805 & ~w12806;
assign w12826 = ~w12819 & ~w12821;
assign w12827 = w12825 & w12826;
assign w12828 = w12824 & w12827;
assign w12829 = w12708 & w12820;
assign w12830 = pi056 & w3321;
assign w12831 = w3369 & w12830;
assign w12832 = pi080 & w3353;
assign w12833 = pi088 & w3402;
assign w12834 = pi040 & w3420;
assign w12835 = pi104 & w4051;
assign w12836 = pi112 & w4071;
assign w12837 = pi096 & w4083;
assign w12838 = ~w12835 & ~w12836;
assign w12839 = ~w12829 & w12838;
assign w12840 = ~w12831 & ~w12832;
assign w12841 = ~w12833 & ~w12834;
assign w12842 = ~w12837 & w12841;
assign w12843 = w12839 & w12840;
assign w12844 = w12842 & w12843;
assign w12845 = w12725 & w12820;
assign w12846 = pi057 & w3321;
assign w12847 = w3369 & w12846;
assign w12848 = pi081 & w3353;
assign w12849 = pi089 & w3402;
assign w12850 = pi041 & w3420;
assign w12851 = pi113 & w4071;
assign w12852 = pi105 & w4051;
assign w12853 = pi097 & w4083;
assign w12854 = ~w12851 & ~w12852;
assign w12855 = ~w12845 & w12854;
assign w12856 = ~w12847 & ~w12848;
assign w12857 = ~w12849 & ~w12850;
assign w12858 = ~w12853 & w12857;
assign w12859 = w12855 & w12856;
assign w12860 = w12858 & w12859;
assign w12861 = pi042 & w3420;
assign w12862 = pi074 & w3387;
assign w12863 = pi098 & w4083;
assign w12864 = pi058 & w4094;
assign w12865 = pi082 & w3353;
assign w12866 = pi114 & w4071;
assign w12867 = pi106 & w4051;
assign w12868 = pi090 & w3402;
assign w12869 = ~w12866 & ~w12867;
assign w12870 = ~w12861 & w12869;
assign w12871 = ~w12862 & ~w12863;
assign w12872 = ~w12864 & ~w12865;
assign w12873 = ~w12868 & w12872;
assign w12874 = w12870 & w12871;
assign w12875 = w12873 & w12874;
assign w12876 = pi059 & w3321;
assign w12877 = w3369 & w12876;
assign w12878 = w12753 & w12820;
assign w12879 = pi091 & w3402;
assign w12880 = pi043 & w3420;
assign w12881 = pi099 & w4083;
assign w12882 = pi115 & w4071;
assign w12883 = pi107 & w4051;
assign w12884 = pi083 & w3353;
assign w12885 = ~w12882 & ~w12883;
assign w12886 = ~w12877 & w12885;
assign w12887 = ~w12878 & ~w12879;
assign w12888 = ~w12880 & ~w12881;
assign w12889 = ~w12884 & w12888;
assign w12890 = w12886 & w12887;
assign w12891 = w12889 & w12890;
assign w12892 = pi060 & w3321;
assign w12893 = w3369 & w12892;
assign w12894 = w12764 & w12820;
assign w12895 = pi092 & w3402;
assign w12896 = pi044 & w3420;
assign w12897 = pi100 & w4083;
assign w12898 = pi108 & w4051;
assign w12899 = pi116 & w4071;
assign w12900 = pi084 & w3353;
assign w12901 = ~w12898 & ~w12899;
assign w12902 = ~w12893 & w12901;
assign w12903 = ~w12894 & ~w12895;
assign w12904 = ~w12896 & ~w12897;
assign w12905 = ~w12900 & w12904;
assign w12906 = w12902 & w12903;
assign w12907 = w12905 & w12906;
assign w12908 = pi061 & w3321;
assign w12909 = w3369 & w12908;
assign w12910 = w12779 & w12820;
assign w12911 = pi101 & w4083;
assign w12912 = pi093 & w3402;
assign w12913 = pi085 & w3353;
assign w12914 = pi109 & w4051;
assign w12915 = pi117 & w4071;
assign w12916 = pi045 & w3420;
assign w12917 = ~w12914 & ~w12915;
assign w12918 = ~w12909 & w12917;
assign w12919 = ~w12910 & ~w12911;
assign w12920 = ~w12912 & ~w12913;
assign w12921 = ~w12916 & w12920;
assign w12922 = w12918 & w12919;
assign w12923 = w12921 & w12922;
assign w12924 = pi078 & w3387;
assign w12925 = pi102 & w4083;
assign w12926 = pi086 & w3353;
assign w12927 = pi094 & w3402;
assign w12928 = pi062 & w4094;
assign w12929 = pi110 & w4051;
assign w12930 = pi118 & w4071;
assign w12931 = pi046 & w3420;
assign w12932 = ~w12929 & ~w12930;
assign w12933 = ~w12924 & w12932;
assign w12934 = ~w12925 & ~w12926;
assign w12935 = ~w12927 & ~w12928;
assign w12936 = ~w12931 & w12935;
assign w12937 = w12933 & w12934;
assign w12938 = w12936 & w12937;
assign w12939 = pi127 & w4742;
assign w12940 = pi055 & w4828;
assign w12941 = pi079 & w4100;
assign w12942 = pi103 & w3948;
assign w12943 = w3977 & w12942;
assign w12944 = w3920 & w12943;
assign w12945 = w4748 & w12944;
assign w12946 = w4755 & w12945;
assign w12947 = w4806 & w12692;
assign w12948 = pi111 & w4783;
assign w12949 = pi095 & w4767;
assign w12950 = w4843 & w4852;
assign w12951 = w12817 & w12950;
assign w12952 = pi119 & w4687;
assign w12953 = w4702 & w12811;
assign w12954 = w4697 & w12953;
assign w12955 = w4694 & w12954;
assign w12956 = ~w12939 & ~w12941;
assign w12957 = ~w12946 & ~w12955;
assign w12958 = w12956 & w12957;
assign w12959 = ~w12940 & ~w12947;
assign w12960 = ~w12948 & ~w12949;
assign w12961 = ~w12951 & ~w12952;
assign w12962 = w12960 & w12961;
assign w12963 = w12958 & w12959;
assign w12964 = w12962 & w12963;
assign w12965 = pi088 & w4705;
assign w12966 = pi120 & w4687;
assign w12967 = pi080 & w4100;
assign w12968 = pi104 & w4757;
assign w12969 = ~w852 & w12950;
assign w12970 = pi040 & w5594;
assign w12971 = w12969 & w12970;
assign w12972 = pi096 & w4767;
assign w12973 = pi112 & w4783;
assign w12974 = w4806 & w12708;
assign w12975 = pi056 & w4828;
assign w12976 = pi128 & w4742;
assign w12977 = ~w12967 & ~w12976;
assign w12978 = ~w12965 & w12977;
assign w12979 = ~w12966 & ~w12968;
assign w12980 = ~w12972 & ~w12973;
assign w12981 = ~w12974 & ~w12975;
assign w12982 = w12980 & w12981;
assign w12983 = w12978 & w12979;
assign w12984 = ~w12971 & w12983;
assign w12985 = w12982 & w12984;
assign w12986 = pi057 & w4828;
assign w12987 = pi097 & w4767;
assign w12988 = pi081 & w4100;
assign w12989 = pi121 & w4687;
assign w12990 = pi041 & w5594;
assign w12991 = w12969 & w12990;
assign w12992 = pi113 & w4783;
assign w12993 = pi105 & w4757;
assign w12994 = w4806 & w12725;
assign w12995 = pi089 & w4705;
assign w12996 = pi129 & w4742;
assign w12997 = ~w12988 & ~w12996;
assign w12998 = ~w12986 & w12997;
assign w12999 = ~w12987 & ~w12989;
assign w13000 = ~w12992 & ~w12993;
assign w13001 = ~w12994 & ~w12995;
assign w13002 = w13000 & w13001;
assign w13003 = w12998 & w12999;
assign w13004 = ~w12991 & w13003;
assign w13005 = w13002 & w13004;
assign w13006 = pi098 & w4767;
assign w13007 = pi090 & w4705;
assign w13008 = pi130 & w4742;
assign w13009 = w4806 & w12736;
assign w13010 = pi042 & w5594;
assign w13011 = w12969 & w13010;
assign w13012 = pi106 & w4757;
assign w13013 = pi122 & w4687;
assign w13014 = pi114 & w4783;
assign w13015 = pi058 & w4828;
assign w13016 = pi082 & w4100;
assign w13017 = ~w13008 & ~w13016;
assign w13018 = ~w13006 & w13017;
assign w13019 = ~w13007 & ~w13009;
assign w13020 = ~w13012 & ~w13013;
assign w13021 = ~w13014 & ~w13015;
assign w13022 = w13020 & w13021;
assign w13023 = w13018 & w13019;
assign w13024 = ~w13011 & w13023;
assign w13025 = w13022 & w13024;
assign w13026 = pi091 & w4705;
assign w13027 = w4806 & w12753;
assign w13028 = pi131 & w4742;
assign w13029 = pi107 & w4757;
assign w13030 = pi043 & w5594;
assign w13031 = w12969 & w13030;
assign w13032 = pi059 & w4828;
assign w13033 = pi115 & w4783;
assign w13034 = pi099 & w4767;
assign w13035 = pi123 & w4687;
assign w13036 = pi083 & w4100;
assign w13037 = ~w13028 & ~w13036;
assign w13038 = ~w13026 & w13037;
assign w13039 = ~w13027 & ~w13029;
assign w13040 = ~w13032 & ~w13033;
assign w13041 = ~w13034 & ~w13035;
assign w13042 = w13040 & w13041;
assign w13043 = w13038 & w13039;
assign w13044 = ~w13031 & w13043;
assign w13045 = w13042 & w13044;
assign w13046 = pi108 & w4757;
assign w13047 = w4806 & w12764;
assign w13048 = pi084 & w4100;
assign w13049 = pi116 & w4783;
assign w13050 = pi044 & w5594;
assign w13051 = w12969 & w13050;
assign w13052 = pi092 & w4705;
assign w13053 = pi100 & w4767;
assign w13054 = pi060 & w4828;
assign w13055 = pi124 & w4687;
assign w13056 = pi132 & w4742;
assign w13057 = ~w13048 & ~w13056;
assign w13058 = ~w13046 & w13057;
assign w13059 = ~w13047 & ~w13049;
assign w13060 = ~w13052 & ~w13053;
assign w13061 = ~w13054 & ~w13055;
assign w13062 = w13060 & w13061;
assign w13063 = w13058 & w13059;
assign w13064 = ~w13051 & w13063;
assign w13065 = w13062 & w13064;
assign w13066 = pi101 & w4767;
assign w13067 = w4806 & w12779;
assign w13068 = pi133 & w4742;
assign w13069 = pi093 & w4705;
assign w13070 = pi045 & w5594;
assign w13071 = w12969 & w13070;
assign w13072 = pi061 & w4828;
assign w13073 = pi109 & w4757;
assign w13074 = pi125 & w4687;
assign w13075 = pi117 & w4783;
assign w13076 = pi085 & w4100;
assign w13077 = ~w13068 & ~w13076;
assign w13078 = ~w13066 & w13077;
assign w13079 = ~w13067 & ~w13069;
assign w13080 = ~w13072 & ~w13073;
assign w13081 = ~w13074 & ~w13075;
assign w13082 = w13080 & w13081;
assign w13083 = w13078 & w13079;
assign w13084 = ~w13071 & w13083;
assign w13085 = w13082 & w13084;
assign w13086 = pi102 & w4767;
assign w13087 = pi110 & w4757;
assign w13088 = pi134 & w4742;
assign w13089 = pi062 & w4828;
assign w13090 = pi046 & w5594;
assign w13091 = w12969 & w13090;
assign w13092 = pi126 & w4687;
assign w13093 = pi094 & w4705;
assign w13094 = w4806 & w12792;
assign w13095 = pi118 & w4783;
assign w13096 = pi086 & w4100;
assign w13097 = ~w13088 & ~w13096;
assign w13098 = ~w13086 & w13097;
assign w13099 = ~w13087 & ~w13089;
assign w13100 = ~w13092 & ~w13093;
assign w13101 = ~w13094 & ~w13095;
assign w13102 = w13100 & w13101;
assign w13103 = w13098 & w13099;
assign w13104 = ~w13091 & w13103;
assign w13105 = w13102 & w13104;
assign w13106 = w5429 & w5442;
assign w13107 = ~w4051 & w12942;
assign w13108 = w13106 & w13107;
assign w13109 = pi087 & w3252;
assign w13110 = w2783 & w13109;
assign w13111 = w2843 & w13110;
assign w13112 = w3169 & w13111;
assign w13113 = ~w2873 & w5527;
assign w13114 = w13112 & w13113;
assign w13115 = w5523 & w13114;
assign w13116 = w5521 & w13115;
assign w13117 = pi119 & w4579;
assign w13118 = w4550 & w13117;
assign w13119 = w4669 & w13118;
assign w13120 = w4522 & w13119;
assign w13121 = w5460 & w13120;
assign w13122 = pi111 & w5422;
assign w13123 = pi127 & w5502;
assign w13124 = pi143 & w5481;
assign w13125 = w1728 & w12613;
assign w13126 = w5584 & w13125;
assign w13127 = w4838 & w12514;
assign w13128 = w5597 & w13127;
assign w13129 = w5610 & w13128;
assign w13130 = pi095 & w5541;
assign w13131 = w911 & w6109;
assign w13132 = ~w906 & w13131;
assign w13133 = w4716 & w13132;
assign w13134 = w5396 & w13133;
assign w13135 = pi071 & ~w2197;
assign w13136 = w1920 & w13135;
assign w13137 = ~w1949 & w13136;
assign w13138 = w5542 & w13137;
assign w13139 = w5562 & w13138;
assign w13140 = ~w13116 & ~w13134;
assign w13141 = ~w13121 & ~w13122;
assign w13142 = ~w13123 & ~w13124;
assign w13143 = ~w13126 & ~w13129;
assign w13144 = ~w13130 & w13143;
assign w13145 = w13141 & w13142;
assign w13146 = ~w13108 & w13140;
assign w13147 = ~w13139 & w13146;
assign w13148 = w13144 & w13145;
assign w13149 = w13147 & w13148;
assign w13150 = pi088 & w5531;
assign w13151 = pi136 & w5407;
assign w13152 = pi128 & w5502;
assign w13153 = pi112 & w5422;
assign w13154 = pi096 & w5541;
assign w13155 = pi144 & w5481;
assign w13156 = pi104 & w5444;
assign w13157 = pi056 & w1756;
assign w13158 = w5584 & w13157;
assign w13159 = pi040 & w5612;
assign w13160 = pi120 & w5461;
assign w13161 = w5563 & w12708;
assign w13162 = ~w13151 & ~w13152;
assign w13163 = ~w13153 & ~w13154;
assign w13164 = ~w13155 & ~w13158;
assign w13165 = w13163 & w13164;
assign w13166 = ~w13150 & w13162;
assign w13167 = ~w13156 & ~w13159;
assign w13168 = ~w13160 & w13167;
assign w13169 = w13165 & w13166;
assign w13170 = ~w13161 & w13169;
assign w13171 = w13168 & w13170;
assign w13172 = pi041 & w5612;
assign w13173 = pi137 & w5407;
assign w13174 = pi113 & w5422;
assign w13175 = pi057 & w5641;
assign w13176 = pi129 & w5502;
assign w13177 = pi097 & w5541;
assign w13178 = pi089 & w5531;
assign w13179 = pi145 & w5481;
assign w13180 = pi121 & w5461;
assign w13181 = pi105 & w5424;
assign w13182 = w13106 & w13181;
assign w13183 = w5563 & w12725;
assign w13184 = ~w13173 & ~w13174;
assign w13185 = ~w13175 & ~w13176;
assign w13186 = ~w13177 & ~w13179;
assign w13187 = w13185 & w13186;
assign w13188 = ~w13172 & w13184;
assign w13189 = ~w13178 & ~w13180;
assign w13190 = ~w13182 & w13189;
assign w13191 = w13187 & w13188;
assign w13192 = ~w13183 & w13191;
assign w13193 = w13190 & w13192;
assign w13194 = pi106 & w5444;
assign w13195 = pi138 & w5407;
assign w13196 = pi098 & w5541;
assign w13197 = pi130 & w5502;
assign w13198 = pi146 & w5481;
assign w13199 = pi058 & w5641;
assign w13200 = pi122 & w5461;
assign w13201 = pi114 & w5422;
assign w13202 = pi042 & w5612;
assign w13203 = pi090 & w5531;
assign w13204 = w5563 & w12736;
assign w13205 = ~w13195 & ~w13196;
assign w13206 = ~w13197 & ~w13198;
assign w13207 = ~w13199 & ~w13201;
assign w13208 = w13206 & w13207;
assign w13209 = ~w13194 & w13205;
assign w13210 = ~w13200 & ~w13202;
assign w13211 = ~w13203 & w13210;
assign w13212 = w13208 & w13209;
assign w13213 = ~w13204 & w13212;
assign w13214 = w13211 & w13213;
assign w13215 = pi043 & w5612;
assign w13216 = pi139 & w5407;
assign w13217 = pi131 & w5502;
assign w13218 = pi147 & w5481;
assign w13219 = pi059 & w1756;
assign w13220 = w5584 & w13219;
assign w13221 = pi099 & w5541;
assign w13222 = pi115 & w5422;
assign w13223 = pi107 & w5444;
assign w13224 = pi091 & w5531;
assign w13225 = pi123 & w5461;
assign w13226 = w5563 & w12753;
assign w13227 = ~w13216 & ~w13217;
assign w13228 = ~w13218 & ~w13220;
assign w13229 = ~w13221 & ~w13222;
assign w13230 = w13228 & w13229;
assign w13231 = ~w13215 & w13227;
assign w13232 = ~w13223 & ~w13224;
assign w13233 = ~w13225 & w13232;
assign w13234 = w13230 & w13231;
assign w13235 = ~w13226 & w13234;
assign w13236 = w13233 & w13235;
assign w13237 = pi108 & w5444;
assign w13238 = pi140 & w5407;
assign w13239 = pi132 & w5502;
assign w13240 = pi060 & w1756;
assign w13241 = w5584 & w13240;
assign w13242 = pi148 & w5481;
assign w13243 = pi100 & w5541;
assign w13244 = pi044 & w5612;
assign w13245 = pi116 & w5422;
assign w13246 = pi124 & w5461;
assign w13247 = pi092 & w5531;
assign w13248 = w5563 & w12764;
assign w13249 = ~w13238 & ~w13239;
assign w13250 = ~w13241 & ~w13242;
assign w13251 = ~w13243 & ~w13245;
assign w13252 = w13250 & w13251;
assign w13253 = ~w13237 & w13249;
assign w13254 = ~w13244 & ~w13246;
assign w13255 = ~w13247 & w13254;
assign w13256 = w13252 & w13253;
assign w13257 = ~w13248 & w13256;
assign w13258 = w13255 & w13257;
assign w13259 = pi125 & w5461;
assign w13260 = pi141 & w5407;
assign w13261 = pi101 & w5541;
assign w13262 = pi061 & w5641;
assign w13263 = pi149 & w5481;
assign w13264 = pi133 & w5502;
assign w13265 = pi093 & w5531;
assign w13266 = pi117 & w5422;
assign w13267 = pi045 & w5612;
assign w13268 = pi109 & w5444;
assign w13269 = w5563 & w12779;
assign w13270 = ~w13260 & ~w13261;
assign w13271 = ~w13262 & ~w13263;
assign w13272 = ~w13264 & ~w13266;
assign w13273 = w13271 & w13272;
assign w13274 = ~w13259 & w13270;
assign w13275 = ~w13265 & ~w13267;
assign w13276 = ~w13268 & w13275;
assign w13277 = w13273 & w13274;
assign w13278 = ~w13269 & w13277;
assign w13279 = w13276 & w13278;
assign w13280 = pi110 & w5444;
assign w13281 = pi142 & w5407;
assign w13282 = pi118 & w5422;
assign w13283 = pi102 & w5541;
assign w13284 = pi150 & w5481;
assign w13285 = pi062 & w5641;
assign w13286 = pi094 & w5531;
assign w13287 = pi134 & w5502;
assign w13288 = pi126 & w5461;
assign w13289 = pi046 & w5612;
assign w13290 = w5563 & w12792;
assign w13291 = ~w13281 & ~w13282;
assign w13292 = ~w13283 & ~w13284;
assign w13293 = ~w13285 & ~w13287;
assign w13294 = w13292 & w13293;
assign w13295 = ~w13280 & w13291;
assign w13296 = ~w13286 & ~w13288;
assign w13297 = ~w13289 & w13296;
assign w13298 = w13294 & w13295;
assign w13299 = ~w13290 & w13298;
assign w13300 = w13297 & w13299;
assign w13301 = pi151 & w6128;
assign w13302 = pi127 & w6308;
assign w13303 = w6335 & w12687;
assign w13304 = w6332 & w13303;
assign w13305 = w6218 & w13114;
assign w13306 = pi143 & w5648;
assign w13307 = pi111 & w6234;
assign w13308 = pi135 & w6170;
assign w13309 = pi095 & w6272;
assign w13310 = w6358 & w12942;
assign w13311 = w6238 & ~w6239;
assign w13312 = w6257 & w13311;
assign w13313 = ~w4831 & w13136;
assign w13314 = w6660 & w13313;
assign w13315 = w13312 & w13314;
assign w13316 = ~w6291 & w13120;
assign w13317 = w6290 & w13316;
assign w13318 = w6287 & w13317;
assign w13319 = pi159 & w6151;
assign w13320 = w6183 & w12514;
assign w13321 = ~w6180 & w13320;
assign w13322 = ~w6179 & w13321;
assign w13323 = w6190 & w13322;
assign w13324 = w6178 & w13323;
assign w13325 = ~w13301 & ~w13318;
assign w13326 = ~w13324 & w13325;
assign w13327 = ~w13305 & ~w13306;
assign w13328 = ~w13307 & ~w13308;
assign w13329 = ~w13309 & ~w13310;
assign w13330 = ~w13315 & w13329;
assign w13331 = w13327 & w13328;
assign w13332 = ~w13302 & w13326;
assign w13333 = ~w13304 & ~w13319;
assign w13334 = w13332 & w13333;
assign w13335 = w13330 & w13331;
assign w13336 = w13334 & w13335;
assign w13337 = pi104 & w6359;
assign w13338 = pi152 & w6128;
assign w13339 = pi144 & w5648;
assign w13340 = pi096 & w6272;
assign w13341 = pi040 & w6195;
assign w13342 = pi112 & w6234;
assign w13343 = pi136 & w6170;
assign w13344 = w6335 & w12830;
assign w13345 = w6332 & w13344;
assign w13346 = ~w2198 & w13312;
assign w13347 = pi072 & w10045;
assign w13348 = w6660 & w10044;
assign w13349 = w13347 & w13348;
assign w13350 = w13346 & w13349;
assign w13351 = pi120 & w6294;
assign w13352 = pi128 & w6308;
assign w13353 = pi088 & w6219;
assign w13354 = pi160 & w6151;
assign w13355 = ~w13338 & ~w13339;
assign w13356 = ~w13340 & ~w13341;
assign w13357 = ~w13342 & ~w13343;
assign w13358 = ~w13351 & w13357;
assign w13359 = w13355 & w13356;
assign w13360 = ~w13337 & ~w13345;
assign w13361 = ~w13350 & ~w13352;
assign w13362 = ~w13353 & ~w13354;
assign w13363 = w13361 & w13362;
assign w13364 = w13359 & w13360;
assign w13365 = w13358 & w13364;
assign w13366 = w13363 & w13365;
assign w13367 = pi089 & w6219;
assign w13368 = pi073 & w10045;
assign w13369 = w13348 & w13368;
assign w13370 = w13346 & w13369;
assign w13371 = pi145 & w5648;
assign w13372 = pi041 & w6195;
assign w13373 = pi097 & w6272;
assign w13374 = pi137 & w6170;
assign w13375 = pi129 & w6308;
assign w13376 = w6335 & w12846;
assign w13377 = w6332 & w13376;
assign w13378 = pi121 & w6294;
assign w13379 = pi105 & w6359;
assign w13380 = pi161 & w6151;
assign w13381 = pi113 & w6234;
assign w13382 = pi153 & w6128;
assign w13383 = ~w13371 & ~w13382;
assign w13384 = ~w13372 & ~w13373;
assign w13385 = ~w13374 & ~w13378;
assign w13386 = ~w13381 & w13385;
assign w13387 = w13383 & w13384;
assign w13388 = ~w13367 & ~w13370;
assign w13389 = ~w13375 & ~w13377;
assign w13390 = ~w13379 & ~w13380;
assign w13391 = w13389 & w13390;
assign w13392 = w13387 & w13388;
assign w13393 = w13386 & w13392;
assign w13394 = w13391 & w13393;
assign w13395 = pi090 & w6219;
assign w13396 = pi146 & w5648;
assign w13397 = pi042 & w6195;
assign w13398 = pi122 & w6294;
assign w13399 = pi138 & w6170;
assign w13400 = pi130 & w6308;
assign w13401 = pi098 & w6272;
assign w13402 = pi114 & w6234;
assign w13403 = pi106 & w6359;
assign w13404 = pi154 & w6128;
assign w13405 = ~w5592 & w13346;
assign w13406 = w3376 & w10044;
assign w13407 = pi074 & w10045;
assign w13408 = w13406 & w13407;
assign w13409 = w13405 & w13408;
assign w13410 = pi162 & w6151;
assign w13411 = pi058 & w3321;
assign w13412 = w6335 & w13411;
assign w13413 = w6332 & w13412;
assign w13414 = ~w13396 & ~w13404;
assign w13415 = ~w13397 & ~w13398;
assign w13416 = ~w13399 & ~w13401;
assign w13417 = ~w13402 & w13416;
assign w13418 = w13414 & w13415;
assign w13419 = ~w13395 & ~w13400;
assign w13420 = ~w13403 & ~w13410;
assign w13421 = ~w13413 & w13420;
assign w13422 = w13418 & w13419;
assign w13423 = ~w13409 & w13417;
assign w13424 = w13422 & w13423;
assign w13425 = w13421 & w13424;
assign w13426 = pi075 & w10045;
assign w13427 = w13406 & w13426;
assign w13428 = w13405 & w13427;
assign w13429 = pi155 & w6128;
assign w13430 = pi099 & w6272;
assign w13431 = pi131 & w6308;
assign w13432 = pi123 & w6294;
assign w13433 = pi043 & w6195;
assign w13434 = pi115 & w6234;
assign w13435 = pi139 & w6170;
assign w13436 = w6335 & w12876;
assign w13437 = w6332 & w13436;
assign w13438 = pi147 & w5648;
assign w13439 = pi091 & w6219;
assign w13440 = pi107 & w6359;
assign w13441 = pi163 & w6151;
assign w13442 = ~w13429 & ~w13430;
assign w13443 = ~w13432 & ~w13433;
assign w13444 = ~w13434 & ~w13435;
assign w13445 = ~w13438 & w13444;
assign w13446 = w13442 & w13443;
assign w13447 = ~w13431 & ~w13437;
assign w13448 = ~w13439 & ~w13440;
assign w13449 = ~w13441 & w13448;
assign w13450 = w13446 & w13447;
assign w13451 = ~w13428 & w13445;
assign w13452 = w13450 & w13451;
assign w13453 = w13449 & w13452;
assign w13454 = pi076 & w10045;
assign w13455 = w13406 & w13454;
assign w13456 = w13405 & w13455;
assign w13457 = pi156 & w6128;
assign w13458 = pi100 & w6272;
assign w13459 = pi092 & w6219;
assign w13460 = pi148 & w5648;
assign w13461 = pi140 & w6170;
assign w13462 = pi116 & w6234;
assign w13463 = pi044 & w6195;
assign w13464 = pi132 & w6308;
assign w13465 = pi124 & w6294;
assign w13466 = w6335 & w12892;
assign w13467 = w6332 & w13466;
assign w13468 = pi108 & w6359;
assign w13469 = pi164 & w6151;
assign w13470 = ~w13457 & ~w13458;
assign w13471 = ~w13460 & ~w13461;
assign w13472 = ~w13462 & ~w13463;
assign w13473 = ~w13465 & w13472;
assign w13474 = w13470 & w13471;
assign w13475 = ~w13459 & ~w13464;
assign w13476 = ~w13467 & ~w13468;
assign w13477 = ~w13469 & w13476;
assign w13478 = w13474 & w13475;
assign w13479 = ~w13456 & w13473;
assign w13480 = w13478 & w13479;
assign w13481 = w13477 & w13480;
assign w13482 = pi077 & w10045;
assign w13483 = w13406 & w13482;
assign w13484 = w13405 & w13483;
assign w13485 = pi125 & w6294;
assign w13486 = pi141 & w6170;
assign w13487 = pi045 & w6195;
assign w13488 = pi149 & w5648;
assign w13489 = pi093 & w6219;
assign w13490 = pi101 & w6272;
assign w13491 = pi109 & w6359;
assign w13492 = w6335 & w12908;
assign w13493 = w6332 & w13492;
assign w13494 = pi133 & w6308;
assign w13495 = pi165 & w6151;
assign w13496 = pi117 & w6234;
assign w13497 = pi157 & w6128;
assign w13498 = ~w13485 & ~w13497;
assign w13499 = ~w13486 & ~w13487;
assign w13500 = ~w13488 & ~w13490;
assign w13501 = ~w13496 & w13500;
assign w13502 = w13498 & w13499;
assign w13503 = ~w13489 & ~w13491;
assign w13504 = ~w13493 & ~w13494;
assign w13505 = ~w13495 & w13504;
assign w13506 = w13502 & w13503;
assign w13507 = ~w13484 & w13501;
assign w13508 = w13506 & w13507;
assign w13509 = w13505 & w13508;
assign w13510 = pi078 & w10045;
assign w13511 = w13406 & w13510;
assign w13512 = w13405 & w13511;
assign w13513 = pi102 & w6272;
assign w13514 = pi126 & w6294;
assign w13515 = pi046 & w6195;
assign w13516 = pi150 & w5648;
assign w13517 = pi062 & w3321;
assign w13518 = w6335 & w13517;
assign w13519 = w6332 & w13518;
assign w13520 = pi142 & w6170;
assign w13521 = pi094 & w6219;
assign w13522 = pi134 & w6308;
assign w13523 = pi110 & w6359;
assign w13524 = pi166 & w6151;
assign w13525 = pi118 & w6234;
assign w13526 = pi158 & w6128;
assign w13527 = ~w13513 & ~w13526;
assign w13528 = ~w13514 & ~w13515;
assign w13529 = ~w13516 & ~w13520;
assign w13530 = ~w13525 & w13529;
assign w13531 = w13527 & w13528;
assign w13532 = ~w13519 & ~w13521;
assign w13533 = ~w13522 & ~w13523;
assign w13534 = ~w13524 & w13533;
assign w13535 = w13531 & w13532;
assign w13536 = ~w13512 & w13530;
assign w13537 = w13535 & w13536;
assign w13538 = w13534 & w13537;
assign w13539 = pi175 & w7157;
assign w13540 = pi111 & w6533;
assign w13541 = pi159 & w7132;
assign w13542 = w7733 & w13118;
assign w13543 = w7712 & w13542;
assign w13544 = w6517 & w13543;
assign w13545 = pi135 & w6441;
assign w13546 = w7165 & w13112;
assign w13547 = w5527 & ~w6535;
assign w13548 = w6542 & w13547;
assign w13549 = w13546 & w13548;
assign w13550 = w6553 & w13549;
assign w13551 = w7106 & w7109;
assign w13552 = w2104 & w13136;
assign w13553 = w2043 & w13552;
assign w13554 = w3376 & w13553;
assign w13555 = w6620 & w13554;
assign w13556 = w6658 & w13555;
assign w13557 = pi143 & w6462;
assign w13558 = w6653 & w13303;
assign w13559 = w6586 & w7177;
assign w13560 = w6587 & w12513;
assign w13561 = w5595 & w13560;
assign w13562 = w6565 & w13561;
assign w13563 = w13559 & w13562;
assign w13564 = pi127 & w6685;
assign w13565 = pi151 & w5888;
assign w13566 = w5948 & w13565;
assign w13567 = w6068 & w13566;
assign w13568 = ~w6128 & w13567;
assign w13569 = w6416 & w13568;
assign w13570 = w6485 & w6492;
assign w13571 = w13107 & w13570;
assign w13572 = ~w13540 & ~w13551;
assign w13573 = ~w13541 & ~w13544;
assign w13574 = ~w13545 & ~w13550;
assign w13575 = ~w13556 & ~w13557;
assign w13576 = ~w13558 & ~w13564;
assign w13577 = ~w13569 & w13576;
assign w13578 = w13574 & w13575;
assign w13579 = w13572 & w13573;
assign w13580 = ~w13539 & ~w13571;
assign w13581 = w13579 & w13580;
assign w13582 = w13577 & w13578;
assign w13583 = ~w13563 & w13582;
assign w13584 = w13581 & w13583;
assign w13585 = pi152 & w6375;
assign w13586 = w6416 & w13585;
assign w13587 = pi120 & w6523;
assign w13588 = w6653 & w13344;
assign w13589 = pi112 & w6533;
assign w13590 = pi144 & w6462;
assign w13591 = pi136 & w6441;
assign w13592 = pi160 & w7132;
assign w13593 = pi168 & w7113;
assign w13594 = pi128 & ~w6307;
assign w13595 = w6685 & w13594;
assign w13596 = pi104 & w6494;
assign w13597 = w7179 & w13559;
assign w13598 = w12970 & w13597;
assign w13599 = pi176 & w7157;
assign w13600 = pi088 & w6558;
assign w13601 = w6659 & w6661;
assign w13602 = w13349 & w13601;
assign w13603 = ~w13586 & ~w13593;
assign w13604 = ~w13588 & ~w13589;
assign w13605 = ~w13590 & ~w13591;
assign w13606 = ~w13592 & ~w13595;
assign w13607 = ~w13600 & w13606;
assign w13608 = w13604 & w13605;
assign w13609 = ~w13587 & w13603;
assign w13610 = ~w13596 & ~w13599;
assign w13611 = w13609 & w13610;
assign w13612 = w13607 & w13608;
assign w13613 = ~w13602 & w13612;
assign w13614 = ~w13598 & w13611;
assign w13615 = w13613 & w13614;
assign w13616 = pi153 & w6375;
assign w13617 = w6416 & w13616;
assign w13618 = pi177 & w7157;
assign w13619 = pi137 & w6441;
assign w13620 = w6653 & w13376;
assign w13621 = pi129 & ~w6307;
assign w13622 = w6685 & w13621;
assign w13623 = pi145 & w6462;
assign w13624 = pi161 & w7132;
assign w13625 = pi169 & w7113;
assign w13626 = pi113 & w6533;
assign w13627 = pi121 & w6523;
assign w13628 = w12990 & w13597;
assign w13629 = w13181 & w13570;
assign w13630 = pi089 & w6558;
assign w13631 = w13369 & w13601;
assign w13632 = ~w13617 & ~w13625;
assign w13633 = ~w13619 & ~w13620;
assign w13634 = ~w13622 & ~w13623;
assign w13635 = ~w13624 & ~w13626;
assign w13636 = ~w13630 & w13635;
assign w13637 = w13633 & w13634;
assign w13638 = ~w13618 & w13632;
assign w13639 = ~w13627 & ~w13629;
assign w13640 = w13638 & w13639;
assign w13641 = w13636 & w13637;
assign w13642 = ~w13631 & w13641;
assign w13643 = ~w13628 & w13640;
assign w13644 = w13642 & w13643;
assign w13645 = pi090 & w6558;
assign w13646 = pi178 & w7157;
assign w13647 = pi138 & w6441;
assign w13648 = pi170 & w7113;
assign w13649 = pi154 & w6375;
assign w13650 = w6416 & w13649;
assign w13651 = pi130 & w6685;
assign w13652 = pi114 & w6533;
assign w13653 = pi146 & w6462;
assign w13654 = w4669 & w6520;
assign w13655 = ~w4551 & w13654;
assign w13656 = w6517 & w13655;
assign w13657 = pi122 & ~w4580;
assign w13658 = w13656 & w13657;
assign w13659 = w6653 & w13412;
assign w13660 = pi106 & w6494;
assign w13661 = w13010 & w13597;
assign w13662 = ~w5592 & w13601;
assign w13663 = w13408 & w13662;
assign w13664 = pi162 & w7132;
assign w13665 = ~w13645 & ~w13648;
assign w13666 = ~w13647 & ~w13650;
assign w13667 = ~w13651 & ~w13652;
assign w13668 = ~w13653 & ~w13659;
assign w13669 = ~w13664 & w13668;
assign w13670 = w13666 & w13667;
assign w13671 = ~w13646 & w13665;
assign w13672 = ~w13658 & ~w13660;
assign w13673 = w13671 & w13672;
assign w13674 = w13669 & w13670;
assign w13675 = w13673 & w13674;
assign w13676 = ~w13661 & ~w13663;
assign w13677 = w13675 & w13676;
assign w13678 = pi171 & w7113;
assign w13679 = pi091 & w6558;
assign w13680 = pi163 & w7132;
assign w13681 = w6653 & w13436;
assign w13682 = pi139 & w6441;
assign w13683 = pi147 & w6462;
assign w13684 = pi115 & w6533;
assign w13685 = pi155 & w6447;
assign w13686 = pi107 & w6494;
assign w13687 = w13427 & w13662;
assign w13688 = pi179 & w7157;
assign w13689 = w13030 & w13597;
assign w13690 = pi131 & w6685;
assign w13691 = pi123 & ~w4580;
assign w13692 = w13656 & w13691;
assign w13693 = ~w13678 & ~w13679;
assign w13694 = ~w13680 & ~w13681;
assign w13695 = ~w13682 & ~w13683;
assign w13696 = ~w13684 & ~w13685;
assign w13697 = ~w13690 & w13696;
assign w13698 = w13694 & w13695;
assign w13699 = ~w13686 & w13693;
assign w13700 = ~w13688 & ~w13692;
assign w13701 = w13699 & w13700;
assign w13702 = w13697 & w13698;
assign w13703 = w13701 & w13702;
assign w13704 = ~w13687 & ~w13689;
assign w13705 = w13703 & w13704;
assign w13706 = pi132 & ~w6307;
assign w13707 = w6685 & w13706;
assign w13708 = pi180 & w7157;
assign w13709 = pi116 & w6533;
assign w13710 = pi172 & w7113;
assign w13711 = pi156 & w6375;
assign w13712 = w6416 & w13711;
assign w13713 = pi164 & w7132;
assign w13714 = pi092 & w6558;
assign w13715 = pi140 & w6441;
assign w13716 = pi124 & ~w4580;
assign w13717 = w13656 & w13716;
assign w13718 = w6653 & w13466;
assign w13719 = pi108 & w6494;
assign w13720 = w13455 & w13662;
assign w13721 = w13050 & w13597;
assign w13722 = pi148 & w6462;
assign w13723 = ~w13707 & ~w13710;
assign w13724 = ~w13709 & ~w13712;
assign w13725 = ~w13713 & ~w13714;
assign w13726 = ~w13715 & ~w13718;
assign w13727 = ~w13722 & w13726;
assign w13728 = w13724 & w13725;
assign w13729 = ~w13708 & w13723;
assign w13730 = ~w13717 & ~w13719;
assign w13731 = w13729 & w13730;
assign w13732 = w13727 & w13728;
assign w13733 = w13731 & w13732;
assign w13734 = ~w13720 & ~w13721;
assign w13735 = w13733 & w13734;
assign w13736 = pi173 & w7113;
assign w13737 = pi133 & ~w6307;
assign w13738 = w6685 & w13737;
assign w13739 = pi149 & w6462;
assign w13740 = pi093 & w6558;
assign w13741 = w6653 & w13492;
assign w13742 = pi117 & w6533;
assign w13743 = pi157 & w6447;
assign w13744 = pi141 & w6441;
assign w13745 = pi109 & w6494;
assign w13746 = w13483 & w13662;
assign w13747 = pi125 & w6523;
assign w13748 = w13070 & w13597;
assign w13749 = pi165 & w7132;
assign w13750 = pi181 & w7157;
assign w13751 = ~w13736 & ~w13738;
assign w13752 = ~w13739 & ~w13740;
assign w13753 = ~w13741 & ~w13742;
assign w13754 = ~w13743 & ~w13744;
assign w13755 = ~w13749 & w13754;
assign w13756 = w13752 & w13753;
assign w13757 = ~w13745 & w13751;
assign w13758 = ~w13747 & ~w13750;
assign w13759 = w13757 & w13758;
assign w13760 = w13755 & w13756;
assign w13761 = w13759 & w13760;
assign w13762 = ~w13746 & ~w13748;
assign w13763 = w13761 & w13762;
assign w13764 = pi174 & w7113;
assign w13765 = pi134 & ~w6307;
assign w13766 = w6685 & w13765;
assign w13767 = pi118 & w6533;
assign w13768 = pi166 & w7132;
assign w13769 = pi094 & w6558;
assign w13770 = pi142 & w6441;
assign w13771 = pi158 & w6447;
assign w13772 = w6653 & w13518;
assign w13773 = pi126 & ~w4580;
assign w13774 = w13656 & w13773;
assign w13775 = w13511 & w13662;
assign w13776 = pi182 & w7157;
assign w13777 = w13090 & w13597;
assign w13778 = pi150 & w6462;
assign w13779 = pi110 & w6494;
assign w13780 = ~w13764 & ~w13766;
assign w13781 = ~w13767 & ~w13768;
assign w13782 = ~w13769 & ~w13770;
assign w13783 = ~w13771 & ~w13772;
assign w13784 = ~w13778 & w13783;
assign w13785 = w13781 & w13782;
assign w13786 = ~w13774 & w13780;
assign w13787 = ~w13776 & ~w13779;
assign w13788 = w13786 & w13787;
assign w13789 = w13784 & w13785;
assign w13790 = w13788 & w13789;
assign w13791 = ~w13775 & ~w13777;
assign w13792 = w13790 & w13791;
assign w13793 = pi191 & w7648;
assign w13794 = w7730 & w13542;
assign w13795 = pi143 & w7229;
assign w13796 = w7965 & w13562;
assign w13797 = w7885 & w13796;
assign w13798 = pi127 & w7751;
assign w13799 = pi111 & w7795;
assign w13800 = w7930 & w13125;
assign w13801 = pi183 & w7585;
assign w13802 = pi135 & w7696;
assign w13803 = pi167 & w7211;
assign w13804 = w6662 & w13553;
assign w13805 = w7857 & w13804;
assign w13806 = w3566 & w6472;
assign w13807 = ~w6494 & w13806;
assign w13808 = w7778 & w13807;
assign w13809 = w7775 & w13808;
assign w13810 = w13107 & w13809;
assign w13811 = pi175 & w7624;
assign w13812 = pi159 & w7603;
assign w13813 = w7804 & ~w7805;
assign w13814 = w7823 & w13813;
assign w13815 = w5526 & w13546;
assign w13816 = w13814 & w13815;
assign w13817 = w5679 & w5739;
assign w13818 = w13567 & w13817;
assign w13819 = w7633 & w13818;
assign w13820 = w7671 & w13819;
assign w13821 = ~w13795 & ~w13801;
assign w13822 = ~w13797 & ~w13799;
assign w13823 = ~w13811 & ~w13812;
assign w13824 = w13822 & w13823;
assign w13825 = ~w13793 & w13821;
assign w13826 = ~w13794 & ~w13798;
assign w13827 = ~w13800 & ~w13802;
assign w13828 = ~w13803 & ~w13805;
assign w13829 = ~w13810 & ~w13816;
assign w13830 = ~w13820 & w13829;
assign w13831 = w13827 & w13828;
assign w13832 = w13825 & w13826;
assign w13833 = w13824 & w13832;
assign w13834 = w13830 & w13831;
assign w13835 = w13833 & w13834;
assign w13836 = pi184 & w7585;
assign w13837 = pi112 & w7795;
assign w13838 = pi104 & w7783;
assign w13839 = w7930 & w13157;
assign w13840 = pi168 & w7211;
assign w13841 = pi144 & w7229;
assign w13842 = pi192 & w7648;
assign w13843 = pi176 & w7624;
assign w13844 = pi136 & w7696;
assign w13845 = w7750 & w13594;
assign w13846 = w7672 & w13585;
assign w13847 = pi120 & ~w4580;
assign w13848 = w7733 & w13847;
assign w13849 = w7731 & w13848;
assign w13850 = w6566 & w7887;
assign w13851 = w12970 & w13850;
assign w13852 = w2932 & w7806;
assign w13853 = w13814 & w13852;
assign w13854 = pi088 & ~w3225;
assign w13855 = w13853 & w13854;
assign w13856 = w6661 & w10044;
assign w13857 = w7858 & w13856;
assign w13858 = w13347 & w13857;
assign w13859 = pi160 & w7603;
assign w13860 = ~w13836 & ~w13837;
assign w13861 = ~w13841 & ~w13843;
assign w13862 = ~w13845 & ~w13859;
assign w13863 = w13861 & w13862;
assign w13864 = ~w13838 & w13860;
assign w13865 = ~w13839 & ~w13840;
assign w13866 = ~w13842 & ~w13844;
assign w13867 = w13865 & w13866;
assign w13868 = w13863 & w13864;
assign w13869 = ~w13846 & ~w13849;
assign w13870 = ~w13851 & ~w13855;
assign w13871 = w13869 & w13870;
assign w13872 = w13867 & w13868;
assign w13873 = ~w13858 & w13872;
assign w13874 = w13871 & w13873;
assign w13875 = w7750 & w13621;
assign w13876 = pi193 & w7648;
assign w13877 = w13181 & w13809;
assign w13878 = pi169 & w7211;
assign w13879 = pi089 & w7827;
assign w13880 = pi041 & w7967;
assign w13881 = pi177 & w7624;
assign w13882 = pi057 & w1756;
assign w13883 = w7930 & w13882;
assign w13884 = pi161 & w7603;
assign w13885 = pi113 & w7795;
assign w13886 = pi121 & ~w4580;
assign w13887 = w7733 & w13886;
assign w13888 = w7731 & w13887;
assign w13889 = pi145 & w7229;
assign w13890 = w7672 & w13616;
assign w13891 = pi185 & w7585;
assign w13892 = w13368 & w13857;
assign w13893 = pi137 & w7696;
assign w13894 = ~w13875 & ~w13891;
assign w13895 = ~w13881 & ~w13884;
assign w13896 = ~w13885 & ~w13889;
assign w13897 = w13895 & w13896;
assign w13898 = ~w13876 & w13894;
assign w13899 = ~w13877 & ~w13878;
assign w13900 = ~w13879 & ~w13880;
assign w13901 = ~w13883 & ~w13893;
assign w13902 = w13900 & w13901;
assign w13903 = w13898 & w13899;
assign w13904 = ~w13888 & w13897;
assign w13905 = ~w13890 & w13904;
assign w13906 = w13902 & w13903;
assign w13907 = ~w13892 & w13906;
assign w13908 = w13905 & w13907;
assign w13909 = pi130 & w7751;
assign w13910 = pi138 & w7696;
assign w13911 = pi146 & w7229;
assign w13912 = pi090 & w7827;
assign w13913 = pi194 & w7648;
assign w13914 = pi162 & w7603;
assign w13915 = pi178 & w7624;
assign w13916 = pi170 & w7211;
assign w13917 = w7733 & w13657;
assign w13918 = w7731 & w13917;
assign w13919 = pi058 & w1756;
assign w13920 = w7930 & w13919;
assign w13921 = pi114 & w7795;
assign w13922 = pi186 & w7585;
assign w13923 = w7672 & w13649;
assign w13924 = pi106 & w7783;
assign w13925 = pi042 & w7967;
assign w13926 = w13407 & w13857;
assign w13927 = ~w13911 & ~w13922;
assign w13928 = ~w13914 & ~w13915;
assign w13929 = ~w13921 & w13928;
assign w13930 = ~w13909 & w13927;
assign w13931 = ~w13910 & ~w13912;
assign w13932 = ~w13913 & ~w13916;
assign w13933 = ~w13920 & ~w13924;
assign w13934 = ~w13925 & w13933;
assign w13935 = w13931 & w13932;
assign w13936 = w13929 & w13930;
assign w13937 = ~w13918 & ~w13923;
assign w13938 = w13936 & w13937;
assign w13939 = w13934 & w13935;
assign w13940 = ~w13926 & w13939;
assign w13941 = w13938 & w13940;
assign w13942 = pi163 & w7603;
assign w13943 = pi139 & w7696;
assign w13944 = w7930 & w13219;
assign w13945 = pi171 & w7211;
assign w13946 = pi091 & w7827;
assign w13947 = pi107 & w5424;
assign w13948 = w13809 & w13947;
assign w13949 = pi147 & w7229;
assign w13950 = pi131 & w7751;
assign w13951 = pi179 & w7624;
assign w13952 = pi115 & w7795;
assign w13953 = pi155 & w6375;
assign w13954 = w7672 & w13953;
assign w13955 = w13030 & w13850;
assign w13956 = w7733 & w13691;
assign w13957 = w7731 & w13956;
assign w13958 = pi187 & w7585;
assign w13959 = w13426 & w13857;
assign w13960 = pi195 & w7648;
assign w13961 = ~w13942 & ~w13958;
assign w13962 = ~w13949 & ~w13951;
assign w13963 = ~w13952 & w13962;
assign w13964 = ~w13943 & w13961;
assign w13965 = ~w13944 & ~w13945;
assign w13966 = ~w13946 & ~w13948;
assign w13967 = ~w13950 & ~w13960;
assign w13968 = w13966 & w13967;
assign w13969 = w13964 & w13965;
assign w13970 = ~w13954 & w13963;
assign w13971 = ~w13955 & ~w13957;
assign w13972 = w13970 & w13971;
assign w13973 = w13968 & w13969;
assign w13974 = ~w13959 & w13973;
assign w13975 = w13972 & w13974;
assign w13976 = pi188 & w7585;
assign w13977 = pi164 & w7603;
assign w13978 = pi196 & w7648;
assign w13979 = w7930 & w13240;
assign w13980 = pi108 & w7783;
assign w13981 = pi116 & w7795;
assign w13982 = pi172 & w7211;
assign w13983 = pi180 & w7624;
assign w13984 = pi140 & w7696;
assign w13985 = w7750 & w13706;
assign w13986 = w7733 & w13716;
assign w13987 = w7731 & w13986;
assign w13988 = w7672 & w13711;
assign w13989 = w13050 & w13850;
assign w13990 = pi092 & ~w3225;
assign w13991 = w13853 & w13990;
assign w13992 = w13454 & w13857;
assign w13993 = pi148 & w7229;
assign w13994 = ~w13976 & ~w13977;
assign w13995 = ~w13981 & ~w13983;
assign w13996 = ~w13985 & ~w13993;
assign w13997 = w13995 & w13996;
assign w13998 = ~w13978 & w13994;
assign w13999 = ~w13979 & ~w13980;
assign w14000 = ~w13982 & ~w13984;
assign w14001 = w13999 & w14000;
assign w14002 = w13997 & w13998;
assign w14003 = ~w13987 & ~w13988;
assign w14004 = ~w13989 & ~w13991;
assign w14005 = w14003 & w14004;
assign w14006 = w14001 & w14002;
assign w14007 = ~w13992 & w14006;
assign w14008 = w14005 & w14007;
assign w14009 = pi189 & w7585;
assign w14010 = pi117 & w7795;
assign w14011 = pi197 & w7648;
assign w14012 = pi173 & w7211;
assign w14013 = pi141 & w7696;
assign w14014 = pi165 & w7603;
assign w14015 = pi061 & w1756;
assign w14016 = w7930 & w14015;
assign w14017 = pi181 & w7624;
assign w14018 = pi109 & w7783;
assign w14019 = w7750 & w13737;
assign w14020 = w13070 & w13850;
assign w14021 = pi157 & w6375;
assign w14022 = w7672 & w14021;
assign w14023 = pi125 & ~w4580;
assign w14024 = w7733 & w14023;
assign w14025 = w7731 & w14024;
assign w14026 = pi093 & ~w3225;
assign w14027 = w13853 & w14026;
assign w14028 = w13482 & w13857;
assign w14029 = pi149 & w7229;
assign w14030 = ~w14009 & ~w14010;
assign w14031 = ~w14014 & ~w14017;
assign w14032 = ~w14019 & ~w14029;
assign w14033 = w14031 & w14032;
assign w14034 = ~w14011 & w14030;
assign w14035 = ~w14012 & ~w14013;
assign w14036 = ~w14016 & ~w14018;
assign w14037 = w14035 & w14036;
assign w14038 = w14033 & w14034;
assign w14039 = ~w14020 & ~w14022;
assign w14040 = ~w14025 & ~w14027;
assign w14041 = w14039 & w14040;
assign w14042 = w14037 & w14038;
assign w14043 = ~w14028 & w14042;
assign w14044 = w14041 & w14043;
assign w14045 = pi190 & w7585;
assign w14046 = pi118 & w7795;
assign w14047 = pi142 & w7696;
assign w14048 = pi174 & w7211;
assign w14049 = pi110 & w7783;
assign w14050 = pi166 & w7603;
assign w14051 = pi062 & w1756;
assign w14052 = w7930 & w14051;
assign w14053 = pi182 & w7624;
assign w14054 = pi198 & w7648;
assign w14055 = w7750 & w13765;
assign w14056 = w7733 & w13773;
assign w14057 = w7731 & w14056;
assign w14058 = pi158 & w6375;
assign w14059 = w7672 & w14058;
assign w14060 = w13090 & w13850;
assign w14061 = pi094 & ~w3225;
assign w14062 = w13853 & w14061;
assign w14063 = w13510 & w13857;
assign w14064 = pi150 & w7229;
assign w14065 = ~w14045 & ~w14046;
assign w14066 = ~w14050 & ~w14053;
assign w14067 = ~w14055 & ~w14064;
assign w14068 = w14066 & w14067;
assign w14069 = ~w14047 & w14065;
assign w14070 = ~w14048 & ~w14049;
assign w14071 = ~w14052 & ~w14054;
assign w14072 = w14070 & w14071;
assign w14073 = w14068 & w14069;
assign w14074 = ~w14057 & ~w14059;
assign w14075 = ~w14060 & ~w14062;
assign w14076 = w14074 & w14075;
assign w14077 = w14072 & w14073;
assign w14078 = ~w14063 & w14077;
assign w14079 = w14076 & w14078;
assign w14080 = pi207 & w8051;
assign w14081 = pi039 & pi223;
assign w14082 = ~w9598 & w14081;
assign w14083 = w155 & w14082;
assign w14084 = w8967 & w14083;
assign w14085 = w597 & w14084;
assign w14086 = w218 & w14085;
assign w14087 = ~w3346 & w14086;
assign w14088 = w7146 & w14087;
assign w14089 = w8688 & w14088;
assign w14090 = ~w3346 & w8342;
assign w14091 = w13552 & w14090;
assign w14092 = ~w8712 & w8720;
assign w14093 = w14091 & w14092;
assign w14094 = w8711 & w14093;
assign w14095 = w13117 & w13654;
assign w14096 = w8545 & w14095;
assign w14097 = pi159 & w8358;
assign w14098 = w8653 & w13125;
assign w14099 = pi167 & w7990;
assign w14100 = pi191 & w8382;
assign w14101 = pi135 & w4982;
assign w14102 = w8344 & w14101;
assign w14103 = ~w4954 & w5012;
assign w14104 = w5162 & w14103;
assign w14105 = w14102 & w14104;
assign w14106 = w8493 & w14105;
assign w14107 = ~w8435 & w13818;
assign w14108 = ~w8434 & w14107;
assign w14109 = w9010 & w14108;
assign w14110 = w8459 & w14109;
assign w14111 = pi127 & w8512;
assign w14112 = pi143 & w8336;
assign w14113 = w8584 & w13546;
assign w14114 = pi199 & w8319;
assign w14115 = pi183 & w8432;
assign w14116 = pi175 & w8403;
assign w14117 = pi103 & w3858;
assign w14118 = w3918 & w14117;
assign w14119 = w8389 & w14118;
assign w14120 = w3832 & w14119;
assign w14121 = ~w8589 & w8603;
assign w14122 = w14120 & w14121;
assign w14123 = w8618 & w14122;
assign w14124 = ~w14080 & ~w14114;
assign w14125 = ~w14111 & w14124;
assign w14126 = ~w14112 & w14125;
assign w14127 = ~w14089 & ~w14094;
assign w14128 = ~w14096 & ~w14097;
assign w14129 = ~w14098 & ~w14099;
assign w14130 = ~w14100 & ~w14110;
assign w14131 = ~w14113 & ~w14115;
assign w14132 = ~w14116 & ~w14123;
assign w14133 = w14131 & w14132;
assign w14134 = w14129 & w14130;
assign w14135 = w14127 & w14128;
assign w14136 = ~w14106 & w14126;
assign w14137 = w14135 & w14136;
assign w14138 = w14133 & w14134;
assign w14139 = w14137 & w14138;
assign w14140 = pi088 & w8551;
assign w14141 = w8587 & w14140;
assign w14142 = w8653 & w13157;
assign w14143 = pi160 & w8358;
assign w14144 = pi208 & w8051;
assign w14145 = pi128 & w8512;
assign w14146 = pi200 & w8319;
assign w14147 = pi144 & w8336;
assign w14148 = pi072 & w8723;
assign w14149 = pi192 & w8382;
assign w14150 = pi184 & w8432;
assign w14151 = pi176 & w8403;
assign w14152 = pi104 & w8621;
assign w14153 = w8460 & w13585;
assign w14154 = w6566 & w8688;
assign w14155 = w12970 & w14154;
assign w14156 = pi168 & w7990;
assign w14157 = w8546 & w13848;
assign w14158 = pi136 & w8463;
assign w14159 = w8493 & w14158;
assign w14160 = ~w14144 & ~w14146;
assign w14161 = ~w14145 & w14160;
assign w14162 = ~w14147 & w14161;
assign w14163 = ~w14142 & ~w14143;
assign w14164 = ~w14148 & ~w14149;
assign w14165 = ~w14150 & ~w14151;
assign w14166 = ~w14152 & ~w14156;
assign w14167 = w14165 & w14166;
assign w14168 = w14163 & w14164;
assign w14169 = ~w14141 & w14162;
assign w14170 = ~w14153 & ~w14155;
assign w14171 = ~w14157 & ~w14159;
assign w14172 = w14170 & w14171;
assign w14173 = w14168 & w14169;
assign w14174 = w14167 & w14173;
assign w14175 = w14172 & w14174;
assign w14176 = pi201 & w8319;
assign w14177 = w8653 & w13882;
assign w14178 = pi209 & w8051;
assign w14179 = pi041 & w9022;
assign w14180 = pi161 & w8358;
assign w14181 = pi193 & w8382;
assign w14182 = pi129 & w8512;
assign w14183 = pi105 & w8621;
assign w14184 = w8460 & w13616;
assign w14185 = pi185 & w8432;
assign w14186 = pi073 & w8723;
assign w14187 = pi089 & w8551;
assign w14188 = w8587 & w14187;
assign w14189 = w8546 & w13887;
assign w14190 = pi137 & w8463;
assign w14191 = w8493 & w14190;
assign w14192 = pi169 & w7990;
assign w14193 = pi177 & w8403;
assign w14194 = pi145 & w8336;
assign w14195 = ~w14176 & ~w14178;
assign w14196 = ~w14182 & w14195;
assign w14197 = ~w14194 & w14196;
assign w14198 = ~w14177 & ~w14179;
assign w14199 = ~w14180 & ~w14181;
assign w14200 = ~w14183 & ~w14185;
assign w14201 = ~w14186 & ~w14192;
assign w14202 = ~w14193 & w14201;
assign w14203 = w14199 & w14200;
assign w14204 = w14197 & w14198;
assign w14205 = ~w14184 & ~w14188;
assign w14206 = ~w14189 & ~w14191;
assign w14207 = w14205 & w14206;
assign w14208 = w14203 & w14204;
assign w14209 = w14202 & w14208;
assign w14210 = w14207 & w14209;
assign w14211 = pi202 & w8319;
assign w14212 = pi074 & w8723;
assign w14213 = pi210 & w8051;
assign w14214 = pi186 & w8432;
assign w14215 = pi178 & w8403;
assign w14216 = pi042 & w9022;
assign w14217 = pi130 & w8512;
assign w14218 = pi058 & w9046;
assign w14219 = pi138 & w8463;
assign w14220 = w8493 & w14219;
assign w14221 = pi170 & w7990;
assign w14222 = pi106 & w8621;
assign w14223 = pi090 & w8551;
assign w14224 = w8587 & w14223;
assign w14225 = w8460 & w13649;
assign w14226 = w8546 & w13917;
assign w14227 = pi194 & w8382;
assign w14228 = pi162 & w8358;
assign w14229 = pi146 & w8336;
assign w14230 = ~w14211 & ~w14213;
assign w14231 = ~w14217 & w14230;
assign w14232 = ~w14229 & w14231;
assign w14233 = ~w14212 & ~w14214;
assign w14234 = ~w14215 & ~w14216;
assign w14235 = ~w14221 & ~w14222;
assign w14236 = ~w14227 & ~w14228;
assign w14237 = w14235 & w14236;
assign w14238 = w14233 & w14234;
assign w14239 = ~w14218 & w14232;
assign w14240 = ~w14220 & ~w14224;
assign w14241 = ~w14225 & ~w14226;
assign w14242 = w14240 & w14241;
assign w14243 = w14238 & w14239;
assign w14244 = w14237 & w14243;
assign w14245 = w14242 & w14244;
assign w14246 = w8546 & w13956;
assign w14247 = w8653 & w13219;
assign w14248 = pi195 & w8382;
assign w14249 = pi211 & w8051;
assign w14250 = pi147 & w8336;
assign w14251 = pi203 & w8319;
assign w14252 = pi131 & w8512;
assign w14253 = pi171 & w7990;
assign w14254 = pi187 & w8432;
assign w14255 = pi179 & w8403;
assign w14256 = pi107 & w8621;
assign w14257 = pi075 & w8723;
assign w14258 = pi139 & w8463;
assign w14259 = w8493 & w14258;
assign w14260 = w8460 & w13953;
assign w14261 = pi163 & w8358;
assign w14262 = w13030 & w14154;
assign w14263 = pi091 & w8551;
assign w14264 = w8587 & w14263;
assign w14265 = ~w14249 & ~w14251;
assign w14266 = ~w14250 & w14265;
assign w14267 = ~w14252 & w14266;
assign w14268 = ~w14247 & ~w14248;
assign w14269 = ~w14253 & ~w14254;
assign w14270 = ~w14255 & ~w14256;
assign w14271 = ~w14257 & ~w14261;
assign w14272 = w14270 & w14271;
assign w14273 = w14268 & w14269;
assign w14274 = ~w14246 & w14267;
assign w14275 = ~w14259 & ~w14260;
assign w14276 = ~w14262 & ~w14264;
assign w14277 = w14275 & w14276;
assign w14278 = w14273 & w14274;
assign w14279 = w14272 & w14278;
assign w14280 = w14277 & w14279;
assign w14281 = pi140 & w8463;
assign w14282 = w8493 & w14281;
assign w14283 = w8653 & w13240;
assign w14284 = pi196 & w8382;
assign w14285 = pi204 & w8319;
assign w14286 = pi148 & w8336;
assign w14287 = pi212 & w8051;
assign w14288 = pi132 & w8512;
assign w14289 = pi188 & w8432;
assign w14290 = pi076 & w8723;
assign w14291 = pi164 & w8358;
assign w14292 = pi180 & w8403;
assign w14293 = pi108 & w8621;
assign w14294 = w8460 & w13711;
assign w14295 = w13050 & w14154;
assign w14296 = pi172 & w7990;
assign w14297 = w8546 & w13986;
assign w14298 = pi092 & w8551;
assign w14299 = w8587 & w14298;
assign w14300 = ~w14285 & ~w14287;
assign w14301 = ~w14286 & w14300;
assign w14302 = ~w14288 & w14301;
assign w14303 = ~w14283 & ~w14284;
assign w14304 = ~w14289 & ~w14290;
assign w14305 = ~w14291 & ~w14292;
assign w14306 = ~w14293 & ~w14296;
assign w14307 = w14305 & w14306;
assign w14308 = w14303 & w14304;
assign w14309 = ~w14282 & w14302;
assign w14310 = ~w14294 & ~w14295;
assign w14311 = ~w14297 & ~w14299;
assign w14312 = w14310 & w14311;
assign w14313 = w14308 & w14309;
assign w14314 = w14307 & w14313;
assign w14315 = w14312 & w14314;
assign w14316 = pi141 & w8463;
assign w14317 = w8493 & w14316;
assign w14318 = w8653 & w14015;
assign w14319 = pi189 & w8432;
assign w14320 = pi205 & w8319;
assign w14321 = pi149 & w8336;
assign w14322 = pi213 & w8051;
assign w14323 = pi133 & w8512;
assign w14324 = pi197 & w8382;
assign w14325 = pi181 & w8403;
assign w14326 = pi173 & w7990;
assign w14327 = pi077 & w8723;
assign w14328 = pi165 & w8358;
assign w14329 = w8460 & w14021;
assign w14330 = w8546 & w14024;
assign w14331 = pi109 & w8621;
assign w14332 = w13070 & w14154;
assign w14333 = pi093 & w8551;
assign w14334 = w8587 & w14333;
assign w14335 = ~w14320 & ~w14322;
assign w14336 = ~w14321 & w14335;
assign w14337 = ~w14323 & w14336;
assign w14338 = ~w14318 & ~w14319;
assign w14339 = ~w14324 & ~w14325;
assign w14340 = ~w14326 & ~w14327;
assign w14341 = ~w14328 & ~w14331;
assign w14342 = w14340 & w14341;
assign w14343 = w14338 & w14339;
assign w14344 = ~w14317 & w14337;
assign w14345 = ~w14329 & ~w14330;
assign w14346 = ~w14332 & ~w14334;
assign w14347 = w14345 & w14346;
assign w14348 = w14343 & w14344;
assign w14349 = w14342 & w14348;
assign w14350 = w14347 & w14349;
assign w14351 = pi142 & w8463;
assign w14352 = w8493 & w14351;
assign w14353 = w8653 & w14051;
assign w14354 = pi190 & w8432;
assign w14355 = pi206 & w8319;
assign w14356 = pi150 & w8336;
assign w14357 = pi214 & w8051;
assign w14358 = pi134 & w8512;
assign w14359 = pi198 & w8382;
assign w14360 = pi166 & w8358;
assign w14361 = pi182 & w8403;
assign w14362 = pi078 & w8723;
assign w14363 = pi174 & w7990;
assign w14364 = w8460 & w14058;
assign w14365 = w8546 & w14056;
assign w14366 = pi110 & w8621;
assign w14367 = w13090 & w14154;
assign w14368 = pi094 & w8551;
assign w14369 = w8587 & w14368;
assign w14370 = ~w14355 & ~w14357;
assign w14371 = ~w14356 & w14370;
assign w14372 = ~w14358 & w14371;
assign w14373 = ~w14353 & ~w14354;
assign w14374 = ~w14359 & ~w14360;
assign w14375 = ~w14361 & ~w14362;
assign w14376 = ~w14363 & ~w14366;
assign w14377 = w14375 & w14376;
assign w14378 = w14373 & w14374;
assign w14379 = ~w14352 & w14372;
assign w14380 = ~w14364 & ~w14365;
assign w14381 = ~w14367 & ~w14369;
assign w14382 = w14380 & w14381;
assign w14383 = w14378 & w14379;
assign w14384 = w14377 & w14383;
assign w14385 = w14382 & w14384;
assign w14386 = w9272 & w14105;
assign w14387 = pi127 & w9325;
assign w14388 = pi191 & w9112;
assign w14389 = w9306 & w14120;
assign w14390 = w9295 & w14389;
assign w14391 = pi143 & w9199;
assign w14392 = pi167 & w9142;
assign w14393 = w9432 & w14091;
assign w14394 = w9414 & w14393;
assign w14395 = w9397 & w13546;
assign w14396 = w10252 & w13117;
assign w14397 = pi199 & w9058;
assign w14398 = pi183 & w9090;
assign w14399 = w9617 & w14081;
assign w14400 = pi215 & w6107;
assign w14401 = w8998 & w14400;
assign w14402 = ~w14399 & ~w14401;
assign w14403 = w8999 & ~w14402;
assign w14404 = pi159 & w9181;
assign w14405 = w9513 & w14085;
assign w14406 = pi175 & w9163;
assign w14407 = pi055 & w9592;
assign w14408 = w9439 & w14407;
assign w14409 = w9447 & w14408;
assign w14410 = w9471 & w14409;
assign w14411 = w9232 & w13568;
assign w14412 = pi207 & w9567;
assign w14413 = ~w14387 & ~w14403;
assign w14414 = ~w14388 & ~w14390;
assign w14415 = ~w14391 & ~w14392;
assign w14416 = ~w14394 & ~w14397;
assign w14417 = ~w14398 & ~w14404;
assign w14418 = ~w14406 & ~w14410;
assign w14419 = w14417 & w14418;
assign w14420 = w14415 & w14416;
assign w14421 = w14413 & w14414;
assign w14422 = ~w14386 & ~w14395;
assign w14423 = ~w14396 & ~w14405;
assign w14424 = ~w14411 & ~w14412;
assign w14425 = w14423 & w14424;
assign w14426 = w14421 & w14422;
assign w14427 = w14419 & w14420;
assign w14428 = w14426 & w14427;
assign w14429 = w14425 & w14428;
assign w14430 = pi072 & w9434;
assign w14431 = pi160 & w9181;
assign w14432 = pi216 & w9005;
assign w14433 = pi192 & w9112;
assign w14434 = pi144 & w9199;
assign w14435 = pi224 & w9621;
assign w14436 = pi168 & w9142;
assign w14437 = w10252 & w13847;
assign w14438 = pi200 & w9058;
assign w14439 = pi208 & w9567;
assign w14440 = pi176 & w9163;
assign w14441 = w9648 & w12551;
assign w14442 = w9272 & w14158;
assign w14443 = pi184 & w9090;
assign w14444 = pi128 & w9325;
assign w14445 = w9398 & w14140;
assign w14446 = w9232 & w13585;
assign w14447 = pi056 & w9474;
assign w14448 = pi104 & w9308;
assign w14449 = ~w14432 & ~w14435;
assign w14450 = ~w14431 & w14449;
assign w14451 = ~w14433 & ~w14434;
assign w14452 = ~w14436 & ~w14438;
assign w14453 = ~w14440 & ~w14443;
assign w14454 = ~w14444 & w14453;
assign w14455 = w14451 & w14452;
assign w14456 = ~w14430 & w14450;
assign w14457 = ~w14437 & ~w14439;
assign w14458 = ~w14441 & ~w14442;
assign w14459 = ~w14446 & ~w14447;
assign w14460 = ~w14448 & w14459;
assign w14461 = w14457 & w14458;
assign w14462 = w14455 & w14456;
assign w14463 = ~w14445 & w14454;
assign w14464 = w14462 & w14463;
assign w14465 = w14460 & w14461;
assign w14466 = w14464 & w14465;
assign w14467 = pi057 & w9474;
assign w14468 = pi129 & w9325;
assign w14469 = pi225 & w9621;
assign w14470 = pi201 & w9058;
assign w14471 = pi169 & w9142;
assign w14472 = pi217 & w9005;
assign w14473 = pi193 & w9112;
assign w14474 = w9232 & w13616;
assign w14475 = pi145 & w9199;
assign w14476 = pi209 & w9567;
assign w14477 = pi185 & w9090;
assign w14478 = w9272 & w14190;
assign w14479 = w10252 & w13886;
assign w14480 = pi161 & w9181;
assign w14481 = pi177 & w9163;
assign w14482 = w9398 & w14187;
assign w14483 = w9648 & w12559;
assign w14484 = pi105 & w9308;
assign w14485 = pi073 & w9434;
assign w14486 = ~w14469 & ~w14472;
assign w14487 = ~w14468 & w14486;
assign w14488 = ~w14470 & ~w14471;
assign w14489 = ~w14473 & ~w14475;
assign w14490 = ~w14477 & ~w14480;
assign w14491 = ~w14481 & w14490;
assign w14492 = w14488 & w14489;
assign w14493 = ~w14467 & w14487;
assign w14494 = ~w14474 & ~w14476;
assign w14495 = ~w14478 & ~w14479;
assign w14496 = ~w14483 & ~w14484;
assign w14497 = ~w14485 & w14496;
assign w14498 = w14494 & w14495;
assign w14499 = w14492 & w14493;
assign w14500 = ~w14482 & w14491;
assign w14501 = w14499 & w14500;
assign w14502 = w14497 & w14498;
assign w14503 = w14501 & w14502;
assign w14504 = w9648 & w12567;
assign w14505 = pi162 & w9181;
assign w14506 = pi226 & w9621;
assign w14507 = pi178 & w9163;
assign w14508 = pi194 & w9112;
assign w14509 = pi218 & w9005;
assign w14510 = pi202 & w9058;
assign w14511 = w9272 & w14219;
assign w14512 = pi170 & w9142;
assign w14513 = pi074 & w9434;
assign w14514 = pi186 & w9090;
assign w14515 = pi106 & w9308;
assign w14516 = w9232 & w13649;
assign w14517 = pi146 & w9199;
assign w14518 = pi130 & w9325;
assign w14519 = w9398 & w14223;
assign w14520 = pi122 & w9363;
assign w14521 = pi058 & w9474;
assign w14522 = pi210 & w9567;
assign w14523 = ~w14506 & ~w14509;
assign w14524 = ~w14505 & w14523;
assign w14525 = ~w14507 & ~w14508;
assign w14526 = ~w14510 & ~w14512;
assign w14527 = ~w14514 & ~w14517;
assign w14528 = ~w14518 & w14527;
assign w14529 = w14525 & w14526;
assign w14530 = ~w14504 & w14524;
assign w14531 = ~w14511 & ~w14513;
assign w14532 = ~w14515 & ~w14516;
assign w14533 = ~w14520 & ~w14521;
assign w14534 = ~w14522 & w14533;
assign w14535 = w14531 & w14532;
assign w14536 = w14529 & w14530;
assign w14537 = ~w14519 & w14528;
assign w14538 = w14536 & w14537;
assign w14539 = w14534 & w14535;
assign w14540 = w14538 & w14539;
assign w14541 = w9232 & w13953;
assign w14542 = pi179 & w9163;
assign w14543 = pi219 & w9005;
assign w14544 = pi195 & w9112;
assign w14545 = pi147 & w9199;
assign w14546 = pi227 & w9621;
assign w14547 = pi163 & w9181;
assign w14548 = pi059 & w9474;
assign w14549 = pi203 & w9058;
assign w14550 = pi107 & w9308;
assign w14551 = pi171 & w9142;
assign w14552 = w9272 & w14258;
assign w14553 = w10252 & w13691;
assign w14554 = pi187 & w9090;
assign w14555 = pi131 & w9325;
assign w14556 = w9398 & w14263;
assign w14557 = w9648 & w12575;
assign w14558 = pi075 & w9434;
assign w14559 = pi211 & w9567;
assign w14560 = ~w14543 & ~w14546;
assign w14561 = ~w14542 & w14560;
assign w14562 = ~w14544 & ~w14545;
assign w14563 = ~w14547 & ~w14549;
assign w14564 = ~w14551 & ~w14554;
assign w14565 = ~w14555 & w14564;
assign w14566 = w14562 & w14563;
assign w14567 = ~w14541 & w14561;
assign w14568 = ~w14548 & ~w14550;
assign w14569 = ~w14552 & ~w14553;
assign w14570 = ~w14557 & ~w14558;
assign w14571 = ~w14559 & w14570;
assign w14572 = w14568 & w14569;
assign w14573 = w14566 & w14567;
assign w14574 = ~w14556 & w14565;
assign w14575 = w14573 & w14574;
assign w14576 = w14571 & w14572;
assign w14577 = w14575 & w14576;
assign w14578 = w10252 & w13716;
assign w14579 = pi196 & w9112;
assign w14580 = pi228 & w9621;
assign w14581 = pi180 & w9163;
assign w14582 = pi148 & w9199;
assign w14583 = pi220 & w9005;
assign w14584 = pi188 & w9090;
assign w14585 = w9272 & w14281;
assign w14586 = pi172 & w9142;
assign w14587 = pi108 & w9308;
assign w14588 = pi204 & w9058;
assign w14589 = w9648 & w12583;
assign w14590 = w9232 & w13711;
assign w14591 = pi164 & w9181;
assign w14592 = pi132 & w9325;
assign w14593 = w9398 & w14298;
assign w14594 = pi212 & w9567;
assign w14595 = pi076 & w9434;
assign w14596 = pi060 & w9474;
assign w14597 = ~w14580 & ~w14583;
assign w14598 = ~w14579 & w14597;
assign w14599 = ~w14581 & ~w14582;
assign w14600 = ~w14584 & ~w14586;
assign w14601 = ~w14588 & ~w14591;
assign w14602 = ~w14592 & w14601;
assign w14603 = w14599 & w14600;
assign w14604 = ~w14578 & w14598;
assign w14605 = ~w14585 & ~w14587;
assign w14606 = ~w14589 & ~w14590;
assign w14607 = ~w14594 & ~w14595;
assign w14608 = ~w14596 & w14607;
assign w14609 = w14605 & w14606;
assign w14610 = w14603 & w14604;
assign w14611 = ~w14593 & w14602;
assign w14612 = w14610 & w14611;
assign w14613 = w14608 & w14609;
assign w14614 = w14612 & w14613;
assign w14615 = w10252 & w14023;
assign w14616 = pi173 & w9142;
assign w14617 = pi229 & w9621;
assign w14618 = pi165 & w9181;
assign w14619 = pi181 & w9163;
assign w14620 = pi221 & w9005;
assign w14621 = pi205 & w9058;
assign w14622 = w9272 & w14316;
assign w14623 = pi149 & w9199;
assign w14624 = pi061 & w9474;
assign w14625 = pi189 & w9090;
assign w14626 = pi077 & w9434;
assign w14627 = pi213 & w9567;
assign w14628 = pi197 & w9112;
assign w14629 = pi133 & w9325;
assign w14630 = w9398 & w14333;
assign w14631 = w9648 & w12591;
assign w14632 = pi109 & w9308;
assign w14633 = w9232 & w14021;
assign w14634 = ~w14617 & ~w14620;
assign w14635 = ~w14616 & w14634;
assign w14636 = ~w14618 & ~w14619;
assign w14637 = ~w14621 & ~w14623;
assign w14638 = ~w14625 & ~w14628;
assign w14639 = ~w14629 & w14638;
assign w14640 = w14636 & w14637;
assign w14641 = ~w14615 & w14635;
assign w14642 = ~w14622 & ~w14624;
assign w14643 = ~w14626 & ~w14627;
assign w14644 = ~w14631 & ~w14632;
assign w14645 = ~w14633 & w14644;
assign w14646 = w14642 & w14643;
assign w14647 = w14640 & w14641;
assign w14648 = ~w14630 & w14639;
assign w14649 = w14647 & w14648;
assign w14650 = w14645 & w14646;
assign w14651 = w14649 & w14650;
assign w14652 = pi062 & w9474;
assign w14653 = pi206 & w9058;
assign w14654 = pi230 & w9621;
assign w14655 = pi182 & w9163;
assign w14656 = pi198 & w9112;
assign w14657 = pi222 & w9005;
assign w14658 = pi166 & w9181;
assign w14659 = pi110 & w9308;
assign w14660 = pi150 & w9199;
assign w14661 = pi214 & w9567;
assign w14662 = pi174 & w9142;
assign w14663 = w9272 & w14351;
assign w14664 = w9232 & w14058;
assign w14665 = pi134 & w9325;
assign w14666 = pi190 & w9090;
assign w14667 = w9398 & w14368;
assign w14668 = w9648 & w12599;
assign w14669 = pi078 & w9434;
assign w14670 = w10252 & w13773;
assign w14671 = ~w14654 & ~w14657;
assign w14672 = ~w14653 & w14671;
assign w14673 = ~w14655 & ~w14656;
assign w14674 = ~w14658 & ~w14660;
assign w14675 = ~w14662 & ~w14665;
assign w14676 = ~w14666 & w14675;
assign w14677 = w14673 & w14674;
assign w14678 = ~w14652 & w14672;
assign w14679 = ~w14659 & ~w14661;
assign w14680 = ~w14663 & ~w14664;
assign w14681 = ~w14668 & ~w14669;
assign w14682 = ~w14670 & w14681;
assign w14683 = w14679 & w14680;
assign w14684 = w14677 & w14678;
assign w14685 = ~w14667 & w14676;
assign w14686 = w14684 & w14685;
assign w14687 = w14682 & w14683;
assign w14688 = w14686 & w14687;
assign w14689 = pi199 & w9730;
assign w14690 = pi159 & w10203;
assign w14691 = pi127 & w9927;
assign w14692 = pi143 & w9842;
assign w14693 = pi191 & w9752;
assign w14694 = pi239 & w10356;
assign w14695 = pi039 & pi231;
assign w14696 = w10502 & w14695;
assign w14697 = ~w14694 & ~w14696;
assign w14698 = w8999 & ~w14697;
assign w14699 = pi215 & w8775;
assign w14700 = w8954 & w14699;
assign w14701 = w12368 & w14700;
assign w14702 = w9636 & w14701;
assign w14703 = ~w9634 & w14702;
assign w14704 = ~w9633 & w14703;
assign w14705 = w9631 & w14704;
assign w14706 = w9653 & w14705;
assign w14707 = w9665 & w14706;
assign w14708 = pi167 & w6782;
assign w14709 = w6811 & w14708;
assign w14710 = w10175 & w14709;
assign w14711 = w10183 & w14710;
assign w14712 = w10173 & w14711;
assign w14713 = w4953 & w14102;
assign w14714 = w9880 & w14713;
assign w14715 = w9877 & w14714;
assign w14716 = pi119 & w4191;
assign w14717 = w4251 & w14716;
assign w14718 = ~w4687 & w14717;
assign w14719 = w11507 & w14718;
assign w14720 = ~w9901 & w14719;
assign w14721 = w9921 & w14720;
assign w14722 = w9898 & w14721;
assign w14723 = pi223 & w10275;
assign w14724 = ~w7183 & w7888;
assign w14725 = pi039 & ~w562;
assign w14726 = ~w593 & w14725;
assign w14727 = w14724 & w14726;
assign w14728 = w7892 & w9013;
assign w14729 = w14727 & w14728;
assign w14730 = w9171 & w14729;
assign w14731 = ~w10121 & w14730;
assign w14732 = w10126 & w14731;
assign w14733 = w10120 & w14732;
assign w14734 = w3771 & w14119;
assign w14735 = ~w8621 & w14734;
assign w14736 = w9930 & w14735;
assign w14737 = w9949 & w14736;
assign w14738 = w9963 & w14737;
assign w14739 = pi175 & w10228;
assign w14740 = pi071 & w2101;
assign w14741 = w1918 & w14740;
assign w14742 = w11647 & w14741;
assign w14743 = w14090 & w14742;
assign w14744 = ~w8723 & w14743;
assign w14745 = w1826 & w14744;
assign w14746 = w10043 & w14745;
assign w14747 = w10030 & w14746;
assign w14748 = pi183 & w9785;
assign w14749 = pi207 & w9697;
assign w14750 = w9824 & w13566;
assign w14751 = w9810 & w14750;
assign w14752 = w3137 & w13109;
assign w14753 = w9969 & w14752;
assign w14754 = ~w9968 & w14753;
assign w14755 = w10006 & w14754;
assign w14756 = pi055 & pi271;
assign w14757 = ~w1448 & w14756;
assign w14758 = w1447 & w14757;
assign w14759 = ~w1482 & ~w1545;
assign w14760 = w14758 & w14759;
assign w14761 = ~w1515 & w14760;
assign w14762 = w9436 & w14761;
assign w14763 = ~w9046 & w14762;
assign w14764 = w10059 & w14763;
assign w14765 = w10088 & w14764;
assign w14766 = ~w14691 & ~w14698;
assign w14767 = ~w14692 & w14766;
assign w14768 = ~w14707 & ~w14712;
assign w14769 = w14767 & w14768;
assign w14770 = ~w14689 & ~w14690;
assign w14771 = ~w14693 & ~w14715;
assign w14772 = ~w14722 & ~w14733;
assign w14773 = ~w14738 & ~w14739;
assign w14774 = ~w14747 & ~w14748;
assign w14775 = ~w14749 & ~w14751;
assign w14776 = ~w14755 & ~w14765;
assign w14777 = w14775 & w14776;
assign w14778 = w14773 & w14774;
assign w14779 = w14771 & w14772;
assign w14780 = w14769 & w14770;
assign w14781 = ~w14723 & w14780;
assign w14782 = w14778 & w14779;
assign w14783 = w14777 & w14782;
assign w14784 = w14781 & w14783;
assign w14785 = pi088 & w10008;
assign w14786 = pi192 & w9752;
assign w14787 = pi072 & w10052;
assign w14788 = pi120 & w9924;
assign w14789 = pi152 & w9826;
assign w14790 = pi104 & w9966;
assign w14791 = pi168 & w10185;
assign w14792 = pi200 & w9730;
assign w14793 = pi056 & w10090;
assign w14794 = pi184 & w9785;
assign w14795 = pi160 & w10203;
assign w14796 = pi224 & w10275;
assign w14797 = pi208 & w9697;
assign w14798 = pi232 & w10542;
assign w14799 = pi144 & w9842;
assign w14800 = pi240 & w10532;
assign w14801 = pi128 & w9927;
assign w14802 = pi176 & w10228;
assign w14803 = pi216 & w9672;
assign w14804 = pi040 & w10130;
assign w14805 = pi136 & w9882;
assign w14806 = ~w14798 & ~w14800;
assign w14807 = ~w14801 & w14806;
assign w14808 = ~w14799 & w14807;
assign w14809 = ~w14786 & w14808;
assign w14810 = ~w14791 & ~w14792;
assign w14811 = ~w14794 & ~w14795;
assign w14812 = ~w14797 & ~w14802;
assign w14813 = ~w14803 & w14812;
assign w14814 = w14810 & w14811;
assign w14815 = ~w14785 & w14809;
assign w14816 = ~w14787 & ~w14788;
assign w14817 = ~w14789 & ~w14790;
assign w14818 = ~w14793 & ~w14796;
assign w14819 = ~w14804 & ~w14805;
assign w14820 = w14818 & w14819;
assign w14821 = w14816 & w14817;
assign w14822 = w14814 & w14815;
assign w14823 = w14813 & w14822;
assign w14824 = w14820 & w14821;
assign w14825 = w14823 & w14824;
assign w14826 = pi073 & w10052;
assign w14827 = pi161 & w10203;
assign w14828 = pi137 & w9882;
assign w14829 = pi225 & w10275;
assign w14830 = pi105 & w9966;
assign w14831 = pi121 & w9924;
assign w14832 = pi217 & w9672;
assign w14833 = pi169 & w10185;
assign w14834 = pi153 & w9826;
assign w14835 = pi185 & w9785;
assign w14836 = pi193 & w9752;
assign w14837 = pi041 & w10130;
assign w14838 = pi201 & w9730;
assign w14839 = pi241 & w10532;
assign w14840 = pi145 & w9842;
assign w14841 = pi233 & w10542;
assign w14842 = pi129 & w9927;
assign w14843 = pi209 & w9697;
assign w14844 = pi177 & w10228;
assign w14845 = pi057 & w10090;
assign w14846 = pi089 & w10008;
assign w14847 = ~w14839 & ~w14841;
assign w14848 = ~w14842 & w14847;
assign w14849 = ~w14840 & w14848;
assign w14850 = ~w14827 & w14849;
assign w14851 = ~w14832 & ~w14833;
assign w14852 = ~w14835 & ~w14836;
assign w14853 = ~w14838 & ~w14843;
assign w14854 = ~w14844 & w14853;
assign w14855 = w14851 & w14852;
assign w14856 = ~w14826 & w14850;
assign w14857 = ~w14828 & ~w14829;
assign w14858 = ~w14830 & ~w14831;
assign w14859 = ~w14834 & ~w14837;
assign w14860 = ~w14845 & ~w14846;
assign w14861 = w14859 & w14860;
assign w14862 = w14857 & w14858;
assign w14863 = w14855 & w14856;
assign w14864 = w14854 & w14863;
assign w14865 = w14861 & w14862;
assign w14866 = w14864 & w14865;
assign w14867 = pi122 & w9924;
assign w14868 = pi170 & w10185;
assign w14869 = pi074 & w10052;
assign w14870 = pi226 & w10275;
assign w14871 = pi106 & w9966;
assign w14872 = pi058 & w10090;
assign w14873 = pi178 & w10228;
assign w14874 = pi210 & w9697;
assign w14875 = pi090 & w10008;
assign w14876 = pi202 & w9730;
assign w14877 = pi186 & w9785;
assign w14878 = pi042 & w10130;
assign w14879 = pi218 & w9672;
assign w14880 = pi234 & w10542;
assign w14881 = pi146 & w9842;
assign w14882 = pi242 & w10532;
assign w14883 = pi130 & w9927;
assign w14884 = pi162 & w10203;
assign w14885 = pi194 & w9752;
assign w14886 = pi138 & w9882;
assign w14887 = pi154 & w9826;
assign w14888 = ~w14880 & ~w14882;
assign w14889 = ~w14883 & w14888;
assign w14890 = ~w14881 & w14889;
assign w14891 = ~w14868 & w14890;
assign w14892 = ~w14873 & ~w14874;
assign w14893 = ~w14876 & ~w14877;
assign w14894 = ~w14879 & ~w14884;
assign w14895 = ~w14885 & w14894;
assign w14896 = w14892 & w14893;
assign w14897 = ~w14867 & w14891;
assign w14898 = ~w14869 & ~w14870;
assign w14899 = ~w14871 & ~w14872;
assign w14900 = ~w14875 & ~w14878;
assign w14901 = ~w14886 & ~w14887;
assign w14902 = w14900 & w14901;
assign w14903 = w14898 & w14899;
assign w14904 = w14896 & w14897;
assign w14905 = w14895 & w14904;
assign w14906 = w14902 & w14903;
assign w14907 = w14905 & w14906;
assign w14908 = pi075 & w10052;
assign w14909 = pi171 & w10185;
assign w14910 = pi139 & w9882;
assign w14911 = pi107 & w9966;
assign w14912 = pi043 & w10130;
assign w14913 = pi059 & w10090;
assign w14914 = pi187 & w9785;
assign w14915 = pi203 & w9730;
assign w14916 = pi155 & w9826;
assign w14917 = pi179 & w10228;
assign w14918 = pi195 & w9752;
assign w14919 = pi091 & w10008;
assign w14920 = pi211 & w9697;
assign w14921 = pi235 & w10542;
assign w14922 = pi147 & w9842;
assign w14923 = pi243 & w10532;
assign w14924 = pi131 & w9927;
assign w14925 = pi219 & w9672;
assign w14926 = pi163 & w10203;
assign w14927 = pi123 & w9924;
assign w14928 = pi227 & w10275;
assign w14929 = ~w14921 & ~w14923;
assign w14930 = ~w14924 & w14929;
assign w14931 = ~w14922 & w14930;
assign w14932 = ~w14909 & w14931;
assign w14933 = ~w14914 & ~w14915;
assign w14934 = ~w14917 & ~w14918;
assign w14935 = ~w14920 & ~w14925;
assign w14936 = ~w14926 & w14935;
assign w14937 = w14933 & w14934;
assign w14938 = ~w14908 & w14932;
assign w14939 = ~w14910 & ~w14911;
assign w14940 = ~w14912 & ~w14913;
assign w14941 = ~w14916 & ~w14919;
assign w14942 = ~w14927 & ~w14928;
assign w14943 = w14941 & w14942;
assign w14944 = w14939 & w14940;
assign w14945 = w14937 & w14938;
assign w14946 = w14936 & w14945;
assign w14947 = w14943 & w14944;
assign w14948 = w14946 & w14947;
assign w14949 = pi156 & w9826;
assign w14950 = pi172 & w10185;
assign w14951 = pi140 & w9882;
assign w14952 = pi228 & w10275;
assign w14953 = pi092 & w10008;
assign w14954 = pi108 & w9966;
assign w14955 = pi220 & w9672;
assign w14956 = pi180 & w10228;
assign w14957 = pi076 & w10052;
assign w14958 = pi164 & w10203;
assign w14959 = pi204 & w9730;
assign w14960 = pi060 & w10090;
assign w14961 = pi196 & w9752;
assign w14962 = pi236 & w10542;
assign w14963 = pi148 & w9842;
assign w14964 = pi244 & w10532;
assign w14965 = pi132 & w9927;
assign w14966 = pi188 & w9785;
assign w14967 = pi212 & w9697;
assign w14968 = pi124 & w9924;
assign w14969 = pi044 & w10130;
assign w14970 = ~w14962 & ~w14964;
assign w14971 = ~w14965 & w14970;
assign w14972 = ~w14963 & w14971;
assign w14973 = ~w14950 & w14972;
assign w14974 = ~w14955 & ~w14956;
assign w14975 = ~w14958 & ~w14959;
assign w14976 = ~w14961 & ~w14966;
assign w14977 = ~w14967 & w14976;
assign w14978 = w14974 & w14975;
assign w14979 = ~w14949 & w14973;
assign w14980 = ~w14951 & ~w14952;
assign w14981 = ~w14953 & ~w14954;
assign w14982 = ~w14957 & ~w14960;
assign w14983 = ~w14968 & ~w14969;
assign w14984 = w14982 & w14983;
assign w14985 = w14980 & w14981;
assign w14986 = w14978 & w14979;
assign w14987 = w14977 & w14986;
assign w14988 = w14984 & w14985;
assign w14989 = w14987 & w14988;
assign w14990 = pi109 & w9966;
assign w14991 = pi189 & w9785;
assign w14992 = pi141 & w9882;
assign w14993 = pi125 & w9924;
assign w14994 = pi077 & w10052;
assign w14995 = pi229 & w10275;
assign w14996 = pi213 & w9697;
assign w14997 = pi173 & w10185;
assign w14998 = pi045 & w10130;
assign w14999 = pi205 & w9730;
assign w15000 = pi181 & w10228;
assign w15001 = pi093 & w10008;
assign w15002 = pi197 & w9752;
assign w15003 = pi245 & w10532;
assign w15004 = pi149 & w9842;
assign w15005 = pi237 & w10542;
assign w15006 = pi133 & w9927;
assign w15007 = pi165 & w10203;
assign w15008 = pi221 & w9672;
assign w15009 = pi061 & w10090;
assign w15010 = pi157 & w9826;
assign w15011 = ~w15003 & ~w15005;
assign w15012 = ~w15006 & w15011;
assign w15013 = ~w15004 & w15012;
assign w15014 = ~w14991 & w15013;
assign w15015 = ~w14996 & ~w14997;
assign w15016 = ~w14999 & ~w15000;
assign w15017 = ~w15002 & ~w15007;
assign w15018 = ~w15008 & w15017;
assign w15019 = w15015 & w15016;
assign w15020 = ~w14990 & w15014;
assign w15021 = ~w14992 & ~w14993;
assign w15022 = ~w14994 & ~w14995;
assign w15023 = ~w14998 & ~w15001;
assign w15024 = ~w15009 & ~w15010;
assign w15025 = w15023 & w15024;
assign w15026 = w15021 & w15022;
assign w15027 = w15019 & w15020;
assign w15028 = w15018 & w15027;
assign w15029 = w15025 & w15026;
assign w15030 = w15028 & w15029;
assign w15031 = pi158 & w9826;
assign w15032 = pi214 & w9697;
assign w15033 = pi078 & w10052;
assign w15034 = pi126 & w9924;
assign w15035 = pi142 & w9882;
assign w15036 = pi230 & w10275;
assign w15037 = pi182 & w10228;
assign w15038 = pi166 & w10203;
assign w15039 = pi046 & w10130;
assign w15040 = pi190 & w9785;
assign w15041 = pi222 & w9672;
assign w15042 = pi062 & w10090;
assign w15043 = pi206 & w9730;
assign w15044 = pi238 & w10542;
assign w15045 = pi150 & w9842;
assign w15046 = pi246 & w10532;
assign w15047 = pi134 & w9927;
assign w15048 = pi198 & w9752;
assign w15049 = pi174 & w10185;
assign w15050 = pi110 & w9966;
assign w15051 = pi094 & w10008;
assign w15052 = ~w15044 & ~w15046;
assign w15053 = ~w15047 & w15052;
assign w15054 = ~w15045 & w15053;
assign w15055 = ~w15032 & w15054;
assign w15056 = ~w15037 & ~w15038;
assign w15057 = ~w15040 & ~w15041;
assign w15058 = ~w15043 & ~w15048;
assign w15059 = ~w15049 & w15058;
assign w15060 = w15056 & w15057;
assign w15061 = ~w15031 & w15055;
assign w15062 = ~w15033 & ~w15034;
assign w15063 = ~w15035 & ~w15036;
assign w15064 = ~w15039 & ~w15042;
assign w15065 = ~w15050 & ~w15051;
assign w15066 = w15064 & w15065;
assign w15067 = w15062 & w15063;
assign w15068 = w15060 & w15061;
assign w15069 = w15059 & w15068;
assign w15070 = w15066 & w15067;
assign w15071 = w15069 & w15070;
assign w15072 = pi207 & w11411;
assign w15073 = pi079 & w10903;
assign w15074 = pi199 & w11366;
assign w15075 = pi191 & w11387;
assign w15076 = pi127 & w11103;
assign w15077 = pi215 & w11440;
assign w15078 = pi175 & w11266;
assign w15079 = pi231 & w10605;
assign w15080 = w10946 & w14727;
assign w15081 = w11067 & w14719;
assign w15082 = w11089 & w15081;
assign w15083 = pi183 & w11246;
assign w15084 = pi095 & w10811;
assign w15085 = pi223 & w10629;
assign w15086 = w10827 & w14753;
assign w15087 = w10852 & w15086;
assign w15088 = w5070 & w14101;
assign w15089 = w11200 & w15088;
assign w15090 = w11195 & w15089;
assign w15091 = w10896 & w14744;
assign w15092 = w10890 & w15091;
assign w15093 = w11118 & w13565;
assign w15094 = w11142 & w15093;
assign w15095 = pi247 & w10804;
assign w15096 = w11020 & w14735;
assign w15097 = w11041 & w15096;
assign w15098 = pi159 & w11323;
assign w15099 = pi143 & w11159;
assign w15100 = pi255 & w10705;
assign w15101 = pi111 & w11048;
assign w15102 = pi239 & w10569;
assign w15103 = ~w10949 & w14763;
assign w15104 = w10964 & w15103;
assign w15105 = w10987 & w15104;
assign w15106 = w11273 & w14710;
assign w15107 = w11304 & w15106;
assign w15108 = ~w15095 & ~w15100;
assign w15109 = ~w15073 & w15108;
assign w15110 = ~w15101 & w15109;
assign w15111 = ~w15084 & w15110;
assign w15112 = ~w15099 & w15111;
assign w15113 = ~w15072 & w15112;
assign w15114 = ~w15074 & ~w15075;
assign w15115 = ~w15076 & ~w15077;
assign w15116 = ~w15078 & ~w15082;
assign w15117 = ~w15083 & ~w15085;
assign w15118 = ~w15087 & ~w15090;
assign w15119 = ~w15092 & ~w15094;
assign w15120 = ~w15097 & ~w15098;
assign w15121 = ~w15102 & ~w15105;
assign w15122 = ~w15107 & w15121;
assign w15123 = w15119 & w15120;
assign w15124 = w15117 & w15118;
assign w15125 = w15115 & w15116;
assign w15126 = w15113 & w15114;
assign w15127 = ~w15079 & ~w15080;
assign w15128 = w15126 & w15127;
assign w15129 = w15124 & w15125;
assign w15130 = w15122 & w15123;
assign w15131 = w15129 & w15130;
assign w15132 = w15128 & w15131;
assign w15133 = pi136 & w11203;
assign w15134 = pi256 & w10705;
assign w15135 = pi088 & w10854;
assign w15136 = pi168 & w11306;
assign w15137 = pi152 & w11144;
assign w15138 = pi072 & w10899;
assign w15139 = pi240 & w10569;
assign w15140 = pi224 & w10629;
assign w15141 = pi144 & w11159;
assign w15142 = pi248 & w10804;
assign w15143 = pi080 & w10903;
assign w15144 = pi128 & w11103;
assign w15145 = pi232 & w10605;
assign w15146 = pi192 & w11387;
assign w15147 = pi160 & w11323;
assign w15148 = pi208 & w11411;
assign w15149 = pi176 & w11266;
assign w15150 = pi112 & w11048;
assign w15151 = pi200 & w11366;
assign w15152 = pi040 & w596;
assign w15153 = w14724 & w15152;
assign w15154 = w10946 & w15153;
assign w15155 = pi184 & w11246;
assign w15156 = pi104 & w11043;
assign w15157 = pi216 & w11440;
assign w15158 = pi096 & w10811;
assign w15159 = pi056 & w10990;
assign w15160 = pi120 & w11091;
assign w15161 = ~w15134 & ~w15142;
assign w15162 = ~w15143 & w15161;
assign w15163 = ~w15150 & w15162;
assign w15164 = ~w15158 & w15163;
assign w15165 = ~w15141 & w15164;
assign w15166 = ~w15139 & w15165;
assign w15167 = ~w15140 & ~w15144;
assign w15168 = ~w15146 & ~w15147;
assign w15169 = ~w15148 & ~w15149;
assign w15170 = ~w15151 & ~w15155;
assign w15171 = ~w15157 & w15170;
assign w15172 = w15168 & w15169;
assign w15173 = w15166 & w15167;
assign w15174 = ~w15133 & ~w15135;
assign w15175 = ~w15136 & ~w15137;
assign w15176 = ~w15138 & ~w15145;
assign w15177 = ~w15154 & ~w15156;
assign w15178 = ~w15159 & ~w15160;
assign w15179 = w15177 & w15178;
assign w15180 = w15175 & w15176;
assign w15181 = w15173 & w15174;
assign w15182 = w15171 & w15172;
assign w15183 = w15181 & w15182;
assign w15184 = w15179 & w15180;
assign w15185 = w15183 & w15184;
assign w15186 = pi137 & w11203;
assign w15187 = pi257 & w10705;
assign w15188 = pi121 & w11091;
assign w15189 = pi089 & w10854;
assign w15190 = pi057 & w10990;
assign w15191 = pi105 & w11043;
assign w15192 = pi201 & w11366;
assign w15193 = pi209 & w11411;
assign w15194 = pi145 & w11159;
assign w15195 = pi249 & w10804;
assign w15196 = pi113 & w11048;
assign w15197 = pi129 & w11103;
assign w15198 = pi153 & w11144;
assign w15199 = pi161 & w11323;
assign w15200 = pi217 & w11440;
assign w15201 = pi225 & w10629;
assign w15202 = pi193 & w11387;
assign w15203 = pi081 & w10903;
assign w15204 = pi241 & w10569;
assign w15205 = pi073 & w10899;
assign w15206 = pi177 & w11266;
assign w15207 = pi233 & w10605;
assign w15208 = pi185 & w11246;
assign w15209 = pi097 & w10811;
assign w15210 = pi041 & w596;
assign w15211 = w14724 & w15210;
assign w15212 = w10946 & w15211;
assign w15213 = pi169 & w11306;
assign w15214 = ~w15187 & ~w15195;
assign w15215 = ~w15196 & w15214;
assign w15216 = ~w15203 & w15215;
assign w15217 = ~w15209 & w15216;
assign w15218 = ~w15194 & w15217;
assign w15219 = ~w15192 & w15218;
assign w15220 = ~w15193 & ~w15197;
assign w15221 = ~w15199 & ~w15200;
assign w15222 = ~w15201 & ~w15202;
assign w15223 = ~w15204 & ~w15206;
assign w15224 = ~w15208 & w15223;
assign w15225 = w15221 & w15222;
assign w15226 = w15219 & w15220;
assign w15227 = ~w15186 & ~w15188;
assign w15228 = ~w15189 & ~w15190;
assign w15229 = ~w15191 & ~w15198;
assign w15230 = ~w15205 & ~w15207;
assign w15231 = ~w15212 & ~w15213;
assign w15232 = w15230 & w15231;
assign w15233 = w15228 & w15229;
assign w15234 = w15226 & w15227;
assign w15235 = w15224 & w15225;
assign w15236 = w15234 & w15235;
assign w15237 = w15232 & w15233;
assign w15238 = w15236 & w15237;
assign w15239 = pi234 & w10605;
assign w15240 = pi250 & w10804;
assign w15241 = pi090 & w10854;
assign w15242 = pi058 & w10990;
assign w15243 = pi106 & w11043;
assign w15244 = pi170 & w11306;
assign w15245 = pi226 & w10629;
assign w15246 = pi194 & w11387;
assign w15247 = pi146 & w11159;
assign w15248 = pi258 & w10705;
assign w15249 = pi114 & w11048;
assign w15250 = pi202 & w11366;
assign w15251 = pi138 & w11203;
assign w15252 = pi242 & w10569;
assign w15253 = pi186 & w11246;
assign w15254 = pi162 & w11323;
assign w15255 = pi178 & w11266;
assign w15256 = pi082 & w10903;
assign w15257 = pi210 & w11411;
assign w15258 = pi122 & w11091;
assign w15259 = pi130 & w11103;
assign w15260 = pi154 & w11144;
assign w15261 = pi218 & w11440;
assign w15262 = pi098 & w10811;
assign w15263 = pi042 & w596;
assign w15264 = w14724 & w15263;
assign w15265 = w10946 & w15264;
assign w15266 = pi074 & w10899;
assign w15267 = ~w15240 & ~w15248;
assign w15268 = ~w15249 & w15267;
assign w15269 = ~w15256 & w15268;
assign w15270 = ~w15262 & w15269;
assign w15271 = ~w15247 & w15270;
assign w15272 = ~w15245 & w15271;
assign w15273 = ~w15246 & ~w15250;
assign w15274 = ~w15252 & ~w15253;
assign w15275 = ~w15254 & ~w15255;
assign w15276 = ~w15257 & ~w15259;
assign w15277 = ~w15261 & w15276;
assign w15278 = w15274 & w15275;
assign w15279 = w15272 & w15273;
assign w15280 = ~w15239 & ~w15241;
assign w15281 = ~w15242 & ~w15243;
assign w15282 = ~w15244 & ~w15251;
assign w15283 = ~w15258 & ~w15260;
assign w15284 = ~w15265 & ~w15266;
assign w15285 = w15283 & w15284;
assign w15286 = w15281 & w15282;
assign w15287 = w15279 & w15280;
assign w15288 = w15277 & w15278;
assign w15289 = w15287 & w15288;
assign w15290 = w15285 & w15286;
assign w15291 = w15289 & w15290;
assign w15292 = pi043 & w596;
assign w15293 = w14724 & w15292;
assign w15294 = w10946 & w15293;
assign w15295 = pi251 & w10804;
assign w15296 = pi075 & w10899;
assign w15297 = pi107 & w11043;
assign w15298 = pi059 & w10990;
assign w15299 = pi171 & w11306;
assign w15300 = pi203 & w11366;
assign w15301 = pi179 & w11266;
assign w15302 = pi147 & w11159;
assign w15303 = pi259 & w10705;
assign w15304 = pi083 & w10903;
assign w15305 = pi187 & w11246;
assign w15306 = pi235 & w10605;
assign w15307 = pi243 & w10569;
assign w15308 = pi219 & w11440;
assign w15309 = pi227 & w10629;
assign w15310 = pi211 & w11411;
assign w15311 = pi115 & w11048;
assign w15312 = pi131 & w11103;
assign w15313 = pi155 & w11144;
assign w15314 = pi163 & w11323;
assign w15315 = pi123 & w11091;
assign w15316 = pi195 & w11387;
assign w15317 = pi099 & w10811;
assign w15318 = pi139 & w11203;
assign w15319 = pi091 & w10854;
assign w15320 = ~w15295 & ~w15303;
assign w15321 = ~w15304 & w15320;
assign w15322 = ~w15311 & w15321;
assign w15323 = ~w15317 & w15322;
assign w15324 = ~w15302 & w15323;
assign w15325 = ~w15300 & w15324;
assign w15326 = ~w15301 & ~w15305;
assign w15327 = ~w15307 & ~w15308;
assign w15328 = ~w15309 & ~w15310;
assign w15329 = ~w15312 & ~w15314;
assign w15330 = ~w15316 & w15329;
assign w15331 = w15327 & w15328;
assign w15332 = w15325 & w15326;
assign w15333 = ~w15294 & ~w15296;
assign w15334 = ~w15297 & ~w15298;
assign w15335 = ~w15299 & ~w15306;
assign w15336 = ~w15313 & ~w15315;
assign w15337 = ~w15318 & ~w15319;
assign w15338 = w15336 & w15337;
assign w15339 = w15334 & w15335;
assign w15340 = w15332 & w15333;
assign w15341 = w15330 & w15331;
assign w15342 = w15340 & w15341;
assign w15343 = w15338 & w15339;
assign w15344 = w15342 & w15343;
assign w15345 = pi124 & w11091;
assign w15346 = pi260 & w10705;
assign w15347 = pi076 & w10899;
assign w15348 = pi156 & w11144;
assign w15349 = pi060 & w10990;
assign w15350 = pi108 & w11043;
assign w15351 = pi132 & w11103;
assign w15352 = pi164 & w11323;
assign w15353 = pi148 & w11159;
assign w15354 = pi252 & w10804;
assign w15355 = pi084 & w10903;
assign w15356 = pi220 & w11440;
assign w15357 = pi172 & w11306;
assign w15358 = pi212 & w11411;
assign w15359 = pi188 & w11246;
assign w15360 = pi244 & w10569;
assign w15361 = pi180 & w11266;
assign w15362 = pi116 & w11048;
assign w15363 = pi228 & w10629;
assign w15364 = pi092 & w10854;
assign w15365 = pi204 & w11366;
assign w15366 = pi140 & w11203;
assign w15367 = pi196 & w11387;
assign w15368 = pi100 & w10811;
assign w15369 = pi044 & w596;
assign w15370 = w14724 & w15369;
assign w15371 = w10946 & w15370;
assign w15372 = pi236 & w10605;
assign w15373 = ~w15346 & ~w15354;
assign w15374 = ~w15355 & w15373;
assign w15375 = ~w15362 & w15374;
assign w15376 = ~w15368 & w15375;
assign w15377 = ~w15353 & w15376;
assign w15378 = ~w15351 & w15377;
assign w15379 = ~w15352 & ~w15356;
assign w15380 = ~w15358 & ~w15359;
assign w15381 = ~w15360 & ~w15361;
assign w15382 = ~w15363 & ~w15365;
assign w15383 = ~w15367 & w15382;
assign w15384 = w15380 & w15381;
assign w15385 = w15378 & w15379;
assign w15386 = ~w15345 & ~w15347;
assign w15387 = ~w15348 & ~w15349;
assign w15388 = ~w15350 & ~w15357;
assign w15389 = ~w15364 & ~w15366;
assign w15390 = ~w15371 & ~w15372;
assign w15391 = w15389 & w15390;
assign w15392 = w15387 & w15388;
assign w15393 = w15385 & w15386;
assign w15394 = w15383 & w15384;
assign w15395 = w15393 & w15394;
assign w15396 = w15391 & w15392;
assign w15397 = w15395 & w15396;
assign w15398 = pi141 & w11203;
assign w15399 = pi253 & w10804;
assign w15400 = pi077 & w10899;
assign w15401 = pi173 & w11306;
assign w15402 = pi061 & w10990;
assign w15403 = pi157 & w11144;
assign w15404 = pi205 & w11366;
assign w15405 = pi197 & w11387;
assign w15406 = pi149 & w11159;
assign w15407 = pi261 & w10705;
assign w15408 = pi117 & w11048;
assign w15409 = pi245 & w10569;
assign w15410 = pi093 & w10854;
assign w15411 = pi229 & w10629;
assign w15412 = pi133 & w11103;
assign w15413 = pi213 & w11411;
assign w15414 = pi181 & w11266;
assign w15415 = pi085 & w10903;
assign w15416 = pi165 & w11323;
assign w15417 = pi125 & w11091;
assign w15418 = pi189 & w11246;
assign w15419 = pi045 & w596;
assign w15420 = w14724 & w15419;
assign w15421 = w10946 & w15420;
assign w15422 = pi221 & w11440;
assign w15423 = pi101 & w10811;
assign w15424 = pi109 & w11043;
assign w15425 = pi237 & w10605;
assign w15426 = ~w15399 & ~w15407;
assign w15427 = ~w15408 & w15426;
assign w15428 = ~w15415 & w15427;
assign w15429 = ~w15423 & w15428;
assign w15430 = ~w15406 & w15429;
assign w15431 = ~w15404 & w15430;
assign w15432 = ~w15405 & ~w15409;
assign w15433 = ~w15411 & ~w15412;
assign w15434 = ~w15413 & ~w15414;
assign w15435 = ~w15416 & ~w15418;
assign w15436 = ~w15422 & w15435;
assign w15437 = w15433 & w15434;
assign w15438 = w15431 & w15432;
assign w15439 = ~w15398 & ~w15400;
assign w15440 = ~w15401 & ~w15402;
assign w15441 = ~w15403 & ~w15410;
assign w15442 = ~w15417 & ~w15421;
assign w15443 = ~w15424 & ~w15425;
assign w15444 = w15442 & w15443;
assign w15445 = w15440 & w15441;
assign w15446 = w15438 & w15439;
assign w15447 = w15436 & w15437;
assign w15448 = w15446 & w15447;
assign w15449 = w15444 & w15445;
assign w15450 = w15448 & w15449;
assign w15451 = pi062 & w10990;
assign w15452 = pi262 & w10705;
assign w15453 = pi094 & w10854;
assign w15454 = pi158 & w11144;
assign w15455 = pi174 & w11306;
assign w15456 = pi078 & w10899;
assign w15457 = pi230 & w10629;
assign w15458 = pi190 & w11246;
assign w15459 = pi150 & w11159;
assign w15460 = pi254 & w10804;
assign w15461 = pi118 & w11048;
assign w15462 = pi214 & w11411;
assign w15463 = pi238 & w10605;
assign w15464 = pi222 & w11440;
assign w15465 = pi182 & w11266;
assign w15466 = pi198 & w11387;
assign w15467 = pi246 & w10569;
assign w15468 = pi086 & w10903;
assign w15469 = pi206 & w11366;
assign w15470 = pi126 & w11091;
assign w15471 = pi166 & w11323;
assign w15472 = pi046 & w596;
assign w15473 = w14724 & w15472;
assign w15474 = w10946 & w15473;
assign w15475 = pi134 & w11103;
assign w15476 = pi102 & w10811;
assign w15477 = pi110 & w11043;
assign w15478 = pi142 & w11203;
assign w15479 = ~w15452 & ~w15460;
assign w15480 = ~w15461 & w15479;
assign w15481 = ~w15468 & w15480;
assign w15482 = ~w15476 & w15481;
assign w15483 = ~w15459 & w15482;
assign w15484 = ~w15457 & w15483;
assign w15485 = ~w15458 & ~w15462;
assign w15486 = ~w15464 & ~w15465;
assign w15487 = ~w15466 & ~w15467;
assign w15488 = ~w15469 & ~w15471;
assign w15489 = ~w15475 & w15488;
assign w15490 = w15486 & w15487;
assign w15491 = w15484 & w15485;
assign w15492 = ~w15451 & ~w15453;
assign w15493 = ~w15454 & ~w15455;
assign w15494 = ~w15456 & ~w15463;
assign w15495 = ~w15470 & ~w15474;
assign w15496 = ~w15477 & ~w15478;
assign w15497 = w15495 & w15496;
assign w15498 = w15493 & w15494;
assign w15499 = w15491 & w15492;
assign w15500 = w15489 & w15490;
assign w15501 = w15499 & w15500;
assign w15502 = w15497 & w15498;
assign w15503 = w15501 & w15502;
assign w15504 = pi239 & w11707;
assign w15505 = pi127 & w12137;
assign w15506 = pi143 & w12251;
assign w15507 = pi159 & w12269;
assign w15508 = w12093 & w14713;
assign w15509 = w12122 & w15508;
assign w15510 = pi223 & w11765;
assign w15511 = pi191 & w12329;
assign w15512 = pi271 & w11635;
assign w15513 = pi263 & w11675;
assign w15514 = pi095 & w12015;
assign w15515 = pi111 & w12006;
assign w15516 = pi255 & w11559;
assign w15517 = pi247 & w11529;
assign w15518 = pi103 & w11996;
assign w15519 = pi199 & w12364;
assign w15520 = w12209 & w13565;
assign w15521 = w12234 & w15520;
assign w15522 = pi231 & w11738;
assign w15523 = w11799 & w11827;
assign w15524 = pi055 & w15523;
assign w15525 = pi071 & w11936;
assign w15526 = pi215 & w12400;
assign w15527 = pi175 & w12481;
assign w15528 = pi079 & w11947;
assign w15529 = w11870 & w11883;
assign w15530 = w14727 & w15529;
assign w15531 = pi167 & w12307;
assign w15532 = pi207 & w12422;
assign w15533 = pi087 & w12072;
assign w15534 = pi119 & w12187;
assign w15535 = pi183 & w12462;
assign w15536 = ~w15512 & ~w15513;
assign w15537 = ~w15505 & w15536;
assign w15538 = ~w15514 & ~w15515;
assign w15539 = ~w15528 & w15538;
assign w15540 = ~w15506 & w15537;
assign w15541 = ~w15507 & ~w15509;
assign w15542 = ~w15521 & w15541;
assign w15543 = w15539 & w15540;
assign w15544 = ~w15504 & ~w15510;
assign w15545 = ~w15511 & ~w15518;
assign w15546 = ~w15519 & ~w15522;
assign w15547 = ~w15524 & ~w15525;
assign w15548 = ~w15526 & ~w15527;
assign w15549 = ~w15530 & ~w15531;
assign w15550 = ~w15532 & ~w15533;
assign w15551 = ~w15534 & ~w15535;
assign w15552 = w15550 & w15551;
assign w15553 = w15548 & w15549;
assign w15554 = w15546 & w15547;
assign w15555 = w15544 & w15545;
assign w15556 = w15542 & w15543;
assign w15557 = ~w15516 & ~w15517;
assign w15558 = w15556 & w15557;
assign w15559 = w15554 & w15555;
assign w15560 = w15552 & w15553;
assign w15561 = w15559 & w15560;
assign w15562 = w15558 & w15561;
assign w15563 = pi056 & w15523;
assign w15564 = pi272 & w11635;
assign w15565 = pi240 & w11707;
assign w15566 = pi200 & w12364;
assign w15567 = pi248 & w11529;
assign w15568 = pi096 & w12015;
assign w15569 = pi080 & w11947;
assign w15570 = pi264 & w11675;
assign w15571 = pi112 & w12006;
assign w15572 = pi104 & w11996;
assign w15573 = pi232 & w11738;
assign w15574 = pi216 & w12400;
assign w15575 = pi088 & w12072;
assign w15576 = w15153 & w15529;
assign w15577 = pi224 & w11765;
assign w15578 = pi120 & w12187;
assign w15579 = pi192 & w12329;
assign w15580 = pi184 & w12462;
assign w15581 = pi072 & w11936;
assign w15582 = pi152 & w12236;
assign w15583 = pi208 & w12422;
assign w15584 = pi176 & w12481;
assign w15585 = pi256 & w11559;
assign w15586 = pi160 & w12269;
assign w15587 = pi136 & w12124;
assign w15588 = pi128 & w12137;
assign w15589 = pi168 & w12307;
assign w15590 = pi144 & w12251;
assign w15591 = ~w15564 & ~w15570;
assign w15592 = ~w15568 & w15591;
assign w15593 = ~w15569 & ~w15571;
assign w15594 = ~w15588 & w15593;
assign w15595 = ~w15586 & w15592;
assign w15596 = ~w15590 & w15595;
assign w15597 = ~w15563 & w15594;
assign w15598 = ~w15565 & ~w15566;
assign w15599 = ~w15572 & ~w15573;
assign w15600 = ~w15574 & ~w15575;
assign w15601 = ~w15576 & ~w15577;
assign w15602 = ~w15578 & ~w15579;
assign w15603 = ~w15580 & ~w15581;
assign w15604 = ~w15582 & ~w15583;
assign w15605 = ~w15584 & ~w15587;
assign w15606 = ~w15589 & w15605;
assign w15607 = w15603 & w15604;
assign w15608 = w15601 & w15602;
assign w15609 = w15599 & w15600;
assign w15610 = w15597 & w15598;
assign w15611 = ~w15567 & w15596;
assign w15612 = ~w15585 & w15611;
assign w15613 = w15609 & w15610;
assign w15614 = w15607 & w15608;
assign w15615 = w15606 & w15614;
assign w15616 = w15612 & w15613;
assign w15617 = w15615 & w15616;
assign w15618 = pi257 & w11559;
assign w15619 = pi105 & w11996;
assign w15620 = pi089 & w12072;
assign w15621 = pi073 & w11936;
assign w15622 = pi185 & w12462;
assign w15623 = pi097 & w12015;
assign w15624 = pi193 & w12329;
assign w15625 = pi201 & w12364;
assign w15626 = pi145 & w12251;
assign w15627 = pi273 & w11635;
assign w15628 = w15211 & w15529;
assign w15629 = pi153 & w12236;
assign w15630 = pi233 & w11738;
assign w15631 = pi249 & w11529;
assign w15632 = pi113 & w12006;
assign w15633 = pi081 & w11947;
assign w15634 = pi265 & w11675;
assign w15635 = pi129 & w12137;
assign w15636 = pi161 & w12269;
assign w15637 = pi121 & w12187;
assign w15638 = pi137 & w12124;
assign w15639 = pi169 & w12307;
assign w15640 = pi209 & w12422;
assign w15641 = pi177 & w12481;
assign w15642 = pi225 & w11765;
assign w15643 = pi217 & w12400;
assign w15644 = pi057 & w15523;
assign w15645 = pi241 & w11707;
assign w15646 = ~w15627 & ~w15634;
assign w15647 = ~w15623 & w15646;
assign w15648 = ~w15632 & ~w15633;
assign w15649 = ~w15635 & w15648;
assign w15650 = ~w15626 & w15647;
assign w15651 = ~w15636 & w15650;
assign w15652 = ~w15619 & w15649;
assign w15653 = ~w15620 & ~w15621;
assign w15654 = ~w15622 & ~w15624;
assign w15655 = ~w15625 & ~w15628;
assign w15656 = ~w15629 & ~w15630;
assign w15657 = ~w15637 & ~w15638;
assign w15658 = ~w15639 & ~w15640;
assign w15659 = ~w15641 & ~w15642;
assign w15660 = ~w15643 & ~w15644;
assign w15661 = ~w15645 & w15660;
assign w15662 = w15658 & w15659;
assign w15663 = w15656 & w15657;
assign w15664 = w15654 & w15655;
assign w15665 = w15652 & w15653;
assign w15666 = ~w15618 & w15651;
assign w15667 = ~w15631 & w15666;
assign w15668 = w15664 & w15665;
assign w15669 = w15662 & w15663;
assign w15670 = w15661 & w15669;
assign w15671 = w15667 & w15668;
assign w15672 = w15670 & w15671;
assign w15673 = pi274 & w11635;
assign w15674 = pi210 & w12422;
assign w15675 = w15264 & w15529;
assign w15676 = pi058 & w15523;
assign w15677 = pi250 & w11529;
assign w15678 = pi130 & w12137;
assign w15679 = pi098 & w12015;
assign w15680 = pi266 & w11675;
assign w15681 = pi114 & w12006;
assign w15682 = pi194 & w12329;
assign w15683 = pi258 & w11559;
assign w15684 = pi234 & w11738;
assign w15685 = pi186 & w12462;
assign w15686 = pi122 & w12187;
assign w15687 = pi170 & w12307;
assign w15688 = pi082 & w11947;
assign w15689 = pi106 & w11996;
assign w15690 = pi162 & w12269;
assign w15691 = pi146 & w12251;
assign w15692 = pi138 & w12124;
assign w15693 = pi090 & w12072;
assign w15694 = pi154 & w12236;
assign w15695 = pi074 & w11936;
assign w15696 = pi226 & w11765;
assign w15697 = pi178 & w12481;
assign w15698 = pi202 & w12364;
assign w15699 = pi218 & w12400;
assign w15700 = pi242 & w11707;
assign w15701 = ~w15673 & ~w15680;
assign w15702 = ~w15678 & w15701;
assign w15703 = ~w15679 & ~w15681;
assign w15704 = ~w15688 & w15703;
assign w15705 = ~w15690 & w15702;
assign w15706 = ~w15691 & w15705;
assign w15707 = ~w15674 & w15704;
assign w15708 = ~w15675 & ~w15676;
assign w15709 = ~w15682 & ~w15684;
assign w15710 = ~w15685 & ~w15686;
assign w15711 = ~w15687 & ~w15689;
assign w15712 = ~w15692 & ~w15693;
assign w15713 = ~w15694 & ~w15695;
assign w15714 = ~w15696 & ~w15697;
assign w15715 = ~w15698 & ~w15699;
assign w15716 = ~w15700 & w15715;
assign w15717 = w15713 & w15714;
assign w15718 = w15711 & w15712;
assign w15719 = w15709 & w15710;
assign w15720 = w15707 & w15708;
assign w15721 = ~w15677 & w15706;
assign w15722 = ~w15683 & w15721;
assign w15723 = w15719 & w15720;
assign w15724 = w15717 & w15718;
assign w15725 = w15716 & w15724;
assign w15726 = w15722 & w15723;
assign w15727 = w15725 & w15726;
assign w15728 = pi275 & w11635;
assign w15729 = pi187 & w12462;
assign w15730 = pi075 & w11936;
assign w15731 = pi059 & w15523;
assign w15732 = pi259 & w11559;
assign w15733 = pi131 & w12137;
assign w15734 = pi099 & w12015;
assign w15735 = pi267 & w11675;
assign w15736 = pi115 & w12006;
assign w15737 = pi195 & w12329;
assign w15738 = pi243 & w11707;
assign w15739 = w15293 & w15529;
assign w15740 = pi235 & w11738;
assign w15741 = pi211 & w12422;
assign w15742 = pi179 & w12481;
assign w15743 = pi083 & w11947;
assign w15744 = pi155 & w12236;
assign w15745 = pi147 & w12251;
assign w15746 = pi163 & w12269;
assign w15747 = pi107 & w11996;
assign w15748 = pi219 & w12400;
assign w15749 = pi203 & w12364;
assign w15750 = pi139 & w12124;
assign w15751 = pi227 & w11765;
assign w15752 = pi171 & w12307;
assign w15753 = pi091 & w12072;
assign w15754 = pi123 & w12187;
assign w15755 = pi251 & w11529;
assign w15756 = ~w15728 & ~w15735;
assign w15757 = ~w15733 & w15756;
assign w15758 = ~w15734 & ~w15736;
assign w15759 = ~w15743 & w15758;
assign w15760 = ~w15745 & w15757;
assign w15761 = ~w15746 & w15760;
assign w15762 = ~w15729 & w15759;
assign w15763 = ~w15730 & ~w15731;
assign w15764 = ~w15737 & ~w15738;
assign w15765 = ~w15739 & ~w15740;
assign w15766 = ~w15741 & ~w15742;
assign w15767 = ~w15744 & ~w15747;
assign w15768 = ~w15748 & ~w15749;
assign w15769 = ~w15750 & ~w15751;
assign w15770 = ~w15752 & ~w15753;
assign w15771 = ~w15754 & w15770;
assign w15772 = w15768 & w15769;
assign w15773 = w15766 & w15767;
assign w15774 = w15764 & w15765;
assign w15775 = w15762 & w15763;
assign w15776 = ~w15732 & w15761;
assign w15777 = ~w15755 & w15776;
assign w15778 = w15774 & w15775;
assign w15779 = w15772 & w15773;
assign w15780 = w15771 & w15779;
assign w15781 = w15777 & w15778;
assign w15782 = w15780 & w15781;
assign w15783 = pi268 & w11675;
assign w15784 = pi244 & w11707;
assign w15785 = pi236 & w11738;
assign w15786 = pi260 & w11559;
assign w15787 = pi132 & w12137;
assign w15788 = pi084 & w11947;
assign w15789 = pi276 & w11635;
assign w15790 = pi116 & w12006;
assign w15791 = pi188 & w12462;
assign w15792 = pi076 & w11936;
assign w15793 = pi172 & w12307;
assign w15794 = pi140 & w12124;
assign w15795 = pi212 & w12422;
assign w15796 = pi220 & w12400;
assign w15797 = pi092 & w12072;
assign w15798 = pi156 & w12236;
assign w15799 = pi148 & w12251;
assign w15800 = pi204 & w12364;
assign w15801 = w15370 & w15529;
assign w15802 = pi100 & w12015;
assign w15803 = pi060 & w15523;
assign w15804 = pi124 & w12187;
assign w15805 = pi252 & w11529;
assign w15806 = pi164 & w12269;
assign w15807 = pi180 & w12481;
assign w15808 = pi108 & w11996;
assign w15809 = pi228 & w11765;
assign w15810 = pi196 & w12329;
assign w15811 = ~w15783 & ~w15789;
assign w15812 = ~w15787 & w15811;
assign w15813 = ~w15788 & ~w15790;
assign w15814 = ~w15802 & w15813;
assign w15815 = ~w15799 & w15812;
assign w15816 = ~w15806 & w15815;
assign w15817 = ~w15784 & w15814;
assign w15818 = ~w15785 & ~w15791;
assign w15819 = ~w15792 & ~w15793;
assign w15820 = ~w15794 & ~w15795;
assign w15821 = ~w15796 & ~w15797;
assign w15822 = ~w15798 & ~w15800;
assign w15823 = ~w15801 & ~w15803;
assign w15824 = ~w15804 & ~w15807;
assign w15825 = ~w15808 & ~w15809;
assign w15826 = ~w15810 & w15825;
assign w15827 = w15823 & w15824;
assign w15828 = w15821 & w15822;
assign w15829 = w15819 & w15820;
assign w15830 = w15817 & w15818;
assign w15831 = ~w15786 & w15816;
assign w15832 = ~w15805 & w15831;
assign w15833 = w15829 & w15830;
assign w15834 = w15827 & w15828;
assign w15835 = w15826 & w15834;
assign w15836 = w15832 & w15833;
assign w15837 = w15835 & w15836;
assign w15838 = pi269 & w11675;
assign w15839 = pi237 & w11738;
assign w15840 = pi093 & w12072;
assign w15841 = pi189 & w12462;
assign w15842 = pi253 & w11529;
assign w15843 = pi101 & w12015;
assign w15844 = pi085 & w11947;
assign w15845 = pi277 & w11635;
assign w15846 = pi133 & w12137;
assign w15847 = pi197 & w12329;
assign w15848 = pi261 & w11559;
assign w15849 = pi141 & w12124;
assign w15850 = pi125 & w12187;
assign w15851 = pi077 & w11936;
assign w15852 = pi173 & w12307;
assign w15853 = pi117 & w12006;
assign w15854 = pi109 & w11996;
assign w15855 = pi149 & w12251;
assign w15856 = pi165 & w12269;
assign w15857 = w15420 & w15529;
assign w15858 = pi213 & w12422;
assign w15859 = pi061 & w15523;
assign w15860 = pi205 & w12364;
assign w15861 = pi229 & w11765;
assign w15862 = pi181 & w12481;
assign w15863 = pi221 & w12400;
assign w15864 = pi157 & w12236;
assign w15865 = pi245 & w11707;
assign w15866 = ~w15838 & ~w15845;
assign w15867 = ~w15843 & w15866;
assign w15868 = ~w15844 & ~w15846;
assign w15869 = ~w15853 & w15868;
assign w15870 = ~w15855 & w15867;
assign w15871 = ~w15856 & w15870;
assign w15872 = ~w15839 & w15869;
assign w15873 = ~w15840 & ~w15841;
assign w15874 = ~w15847 & ~w15849;
assign w15875 = ~w15850 & ~w15851;
assign w15876 = ~w15852 & ~w15854;
assign w15877 = ~w15857 & ~w15858;
assign w15878 = ~w15859 & ~w15860;
assign w15879 = ~w15861 & ~w15862;
assign w15880 = ~w15863 & ~w15864;
assign w15881 = ~w15865 & w15880;
assign w15882 = w15878 & w15879;
assign w15883 = w15876 & w15877;
assign w15884 = w15874 & w15875;
assign w15885 = w15872 & w15873;
assign w15886 = ~w15842 & w15871;
assign w15887 = ~w15848 & w15886;
assign w15888 = w15884 & w15885;
assign w15889 = w15882 & w15883;
assign w15890 = w15881 & w15889;
assign w15891 = w15887 & w15888;
assign w15892 = w15890 & w15891;
assign w15893 = pi190 & w12462;
assign w15894 = pi270 & w11675;
assign w15895 = pi062 & w15523;
assign w15896 = pi078 & w11936;
assign w15897 = pi206 & w12364;
assign w15898 = pi262 & w11559;
assign w15899 = pi102 & w12015;
assign w15900 = pi086 & w11947;
assign w15901 = pi278 & w11635;
assign w15902 = pi118 & w12006;
assign w15903 = pi246 & w11707;
assign w15904 = pi174 & w12307;
assign w15905 = w15473 & w15529;
assign w15906 = pi126 & w12187;
assign w15907 = pi238 & w11738;
assign w15908 = pi134 & w12137;
assign w15909 = pi150 & w12251;
assign w15910 = pi198 & w12329;
assign w15911 = pi166 & w12269;
assign w15912 = pi214 & w12422;
assign w15913 = pi158 & w12236;
assign w15914 = pi094 & w12072;
assign w15915 = pi110 & w11996;
assign w15916 = pi230 & w11765;
assign w15917 = pi142 & w12124;
assign w15918 = pi222 & w12400;
assign w15919 = pi182 & w12481;
assign w15920 = pi254 & w11529;
assign w15921 = ~w15894 & ~w15901;
assign w15922 = ~w15899 & w15921;
assign w15923 = ~w15900 & ~w15902;
assign w15924 = ~w15908 & w15923;
assign w15925 = ~w15909 & w15922;
assign w15926 = ~w15911 & w15925;
assign w15927 = ~w15893 & w15924;
assign w15928 = ~w15895 & ~w15896;
assign w15929 = ~w15897 & ~w15903;
assign w15930 = ~w15904 & ~w15905;
assign w15931 = ~w15906 & ~w15907;
assign w15932 = ~w15910 & ~w15912;
assign w15933 = ~w15913 & ~w15914;
assign w15934 = ~w15915 & ~w15916;
assign w15935 = ~w15917 & ~w15918;
assign w15936 = ~w15919 & w15935;
assign w15937 = w15933 & w15934;
assign w15938 = w15931 & w15932;
assign w15939 = w15929 & w15930;
assign w15940 = w15927 & w15928;
assign w15941 = ~w15898 & w15926;
assign w15942 = ~w15920 & w15941;
assign w15943 = w15939 & w15940;
assign w15944 = w15937 & w15938;
assign w15945 = w15936 & w15944;
assign w15946 = w15942 & w15943;
assign w15947 = w15945 & w15946;
assign w15948 = ~w919 & ~w1759;
assign w15949 = ~w2540 & ~w2552;
assign w15950 = ~w2575 & w15949;
assign w15951 = ~w2552 & ~w2562;
assign w15952 = ~w2590 & ~w3296;
assign w15953 = ~w2635 & ~w3306;
assign w15954 = w15952 & w15953;
assign w15955 = ~w3324 & w15952;
assign w15956 = ~w4051 & ~w4071;
assign w15957 = ~w4083 & w15956;
assign w15958 = ~w3353 & ~w3402;
assign w15959 = ~w3387 & w15958;
assign w15960 = ~w4071 & ~w4094;
assign w15961 = w15958 & w15960;
assign w15962 = ~w4687 & ~w4783;
assign w15963 = ~w4742 & ~w4757;
assign w15964 = ~w4767 & w15963;
assign w15965 = w15962 & w15964;
assign w15966 = ~w4100 & ~w4705;
assign w15967 = ~w4742 & ~w4831;
assign w15968 = w15966 & w15967;
assign w15969 = ~w4828 & w15962;
assign w15970 = w15966 & w15969;
assign w15971 = ~w5407 & ~w5502;
assign w15972 = ~w5422 & ~w5481;
assign w15973 = ~w5461 & w15972;
assign w15974 = ~w5444 & ~w5541;
assign w15975 = w15971 & w15974;
assign w15976 = w15973 & w15975;
assign w15977 = ~w5481 & ~w5592;
assign w15978 = ~w5531 & w15977;
assign w15979 = w15971 & w15978;
assign w15980 = ~w5531 & ~w5641;
assign w15981 = w15973 & w15980;
assign w15982 = ~w6170 & ~w6308;
assign w15983 = ~w5648 & ~w6128;
assign w15984 = ~w6234 & ~w6294;
assign w15985 = w15983 & w15984;
assign w15986 = ~w6272 & ~w6359;
assign w15987 = w15982 & w15986;
assign w15988 = w15985 & w15987;
assign w15989 = ~w6219 & ~w6262;
assign w15990 = w15983 & w15989;
assign w15991 = w15982 & w15990;
assign w15992 = ~w6219 & ~w6381;
assign w15993 = w15985 & w15992;
assign w15994 = ~w7113 & ~w7132;
assign w15995 = ~w7192 & w15994;
assign w15996 = ~w6441 & ~w6685;
assign w15997 = w6463 & ~w6533;
assign w15998 = ~w6523 & w15997;
assign w15999 = ~w6494 & w15996;
assign w16000 = w15998 & w15999;
assign w16001 = w6463 & w6629;
assign w16002 = w15996 & w16001;
assign w16003 = ~w6558 & ~w7172;
assign w16004 = ~w7192 & w16003;
assign w16005 = w15998 & w16004;
assign w16006 = ~w7585 & ~w7624;
assign w16007 = ~w7211 & ~w7603;
assign w16008 = ~w7648 & w16006;
assign w16009 = w16007 & w16008;
assign w16010 = ~w7696 & ~w7751;
assign w16011 = ~w7754 & ~w7795;
assign w16012 = w7702 & ~w7783;
assign w16013 = w16010 & w16011;
assign w16014 = w16012 & w16013;
assign w16015 = w7702 & ~w7827;
assign w16016 = ~w7648 & ~w7899;
assign w16017 = w16010 & w16016;
assign w16018 = w16015 & w16017;
assign w16019 = ~w7960 & w16006;
assign w16020 = w16011 & w16019;
assign w16021 = w16015 & w16020;
assign w16022 = ~w8319 & ~w8382;
assign w16023 = ~w8051 & ~w8403;
assign w16024 = ~w8432 & w16023;
assign w16025 = ~w7990 & ~w8358;
assign w16026 = w16022 & w16025;
assign w16027 = w16024 & w16026;
assign w16028 = w8498 & ~w8512;
assign w16029 = ~w8516 & w16028;
assign w16030 = ~w8548 & ~w8621;
assign w16031 = w16029 & w16030;
assign w16032 = ~w8051 & ~w8658;
assign w16033 = ~w8723 & w16032;
assign w16034 = w16022 & w16033;
assign w16035 = w16029 & w16034;
assign w16036 = w8498 & ~w8658;
assign w16037 = ~w8548 & ~w9046;
assign w16038 = w16036 & w16037;
assign w16039 = w16024 & w16038;
assign w16040 = ~w9090 & ~w9163;
assign w16041 = ~w9005 & ~w9567;
assign w16042 = ~w9058 & ~w9112;
assign w16043 = w16041 & w16042;
assign w16044 = ~w9142 & ~w9621;
assign w16045 = ~w9181 & w16044;
assign w16046 = w16040 & w16045;
assign w16047 = w16043 & w16046;
assign w16048 = w7739 & ~w7740;
assign w16049 = w7747 & w16048;
assign w16050 = w7186 & ~w16049;
assign w16051 = w8468 & ~w16050;
assign w16052 = w8514 & w16051;
assign w16053 = w8492 & w16052;
assign w16054 = ~w9248 & ~w16053;
assign w16055 = w9263 & w16054;
assign w16056 = w9311 & w16055;
assign w16057 = ~w9325 & ~w16056;
assign w16058 = w9240 & w16057;
assign w16059 = ~w9308 & ~w9621;
assign w16060 = ~w9363 & w16059;
assign w16061 = w16058 & w16060;
assign w16062 = ~w9434 & ~w9477;
assign w16063 = w16043 & w16062;
assign w16064 = w16058 & w16063;
assign w16065 = ~w9363 & ~w9474;
assign w16066 = ~w9477 & w16040;
assign w16067 = w16065 & w16066;
assign w16068 = w9240 & w16041;
assign w16069 = w16067 & w16068;
assign w16070 = ~w9785 & ~w10228;
assign w16071 = w10204 & w16070;
assign w16072 = w9754 & w16071;
assign w16073 = ~w10532 & ~w10542;
assign w16074 = ~w10275 & w16073;
assign w16075 = w16072 & w16074;
assign w16076 = ~w9924 & ~w9966;
assign w16077 = ~w9882 & ~w9927;
assign w16078 = w9843 & w16077;
assign w16079 = w16076 & w16078;
assign w16080 = w16072 & ~w16079;
assign w16081 = w16074 & ~w16080;
assign w16082 = ~w10008 & ~w10052;
assign w16083 = w16076 & ~w16082;
assign w16084 = w16078 & ~w16083;
assign w16085 = w16071 & ~w16084;
assign w16086 = w9754 & ~w16085;
assign w16087 = w16074 & ~w16086;
assign w16088 = ~w9924 & ~w10008;
assign w16089 = ~w10090 & w16088;
assign w16090 = w16077 & ~w16089;
assign w16091 = w9843 & ~w16090;
assign w16092 = w10204 & ~w16091;
assign w16093 = w16070 & ~w16092;
assign w16094 = w9753 & ~w16093;
assign w16095 = w9698 & ~w16094;
assign w16096 = ~w10275 & ~w16095;
assign w16097 = ~w10532 & ~w16096;
assign w16098 = w11267 & w11324;
assign w16099 = w11442 & w16098;
assign w16100 = ~w10569 & ~w10804;
assign w16101 = ~w10705 & w16100;
assign w16102 = w10630 & w16101;
assign w16103 = w16099 & w16102;
assign w16104 = w11160 & w11326;
assign w16105 = ~w11048 & ~w11091;
assign w16106 = ~w11043 & w16105;
assign w16107 = ~w10811 & w16104;
assign w16108 = w16106 & w16107;
assign w16109 = w16099 & ~w16108;
assign w16110 = w16102 & ~w16109;
assign w16111 = ~w10854 & ~w10903;
assign w16112 = ~w10899 & w16111;
assign w16113 = w16106 & ~w16112;
assign w16114 = w16104 & ~w16113;
assign w16115 = w16098 & ~w16114;
assign w16116 = w11442 & ~w16115;
assign w16117 = w10631 & ~w16116;
assign w16118 = ~w10705 & ~w16117;
assign w16119 = ~w10990 & w16111;
assign w16120 = ~w11043 & ~w16119;
assign w16121 = w16105 & ~w16120;
assign w16122 = w11326 & ~w16121;
assign w16123 = w11160 & ~w16122;
assign w16124 = w11324 & ~w16123;
assign w16125 = w11267 & ~w16124;
assign w16126 = w11388 & ~w16125;
assign w16127 = w11441 & ~w16126;
assign w16128 = w10630 & ~w16127;
assign w16129 = w16100 & ~w16128;
assign w16130 = ~w12269 & ~w12307;
assign w16131 = w12495 & w16130;
assign w16132 = w12424 & w16131;
assign w16133 = ~w11529 & ~w11707;
assign w16134 = w11766 & w16133;
assign w16135 = ~w11635 & ~w11675;
assign w16136 = ~w11559 & w16135;
assign w16137 = w16134 & w16136;
assign w16138 = w16132 & w16137;
assign w16139 = ~w12006 & ~w12187;
assign w16140 = ~w11996 & w16139;
assign w16141 = w12138 & w12252;
assign w16142 = ~w12015 & w16140;
assign w16143 = w16141 & w16142;
assign w16144 = w16132 & ~w16143;
assign w16145 = w16137 & ~w16144;
assign w16146 = ~w11947 & ~w12072;
assign w16147 = ~w11936 & w16146;
assign w16148 = w16140 & ~w16147;
assign w16149 = (~w16822 & w18153) | (~w16822 & w18154) | (w18153 & w18154);
assign w16150 = w16134 & ~w16149;
assign w16151 = w16136 & ~w16150;
assign w16152 = (~w11996 & ~w16146) | (~w11996 & w16823) | (~w16146 & w16823);
assign w16153 = w16139 & ~w16152;
assign w16154 = w12138 & ~w16153;
assign w16155 = w12252 & w12495;
assign w16156 = ~w16154 & w16155;
assign w16157 = w11559 & ~w11635;
assign w16158 = w12495 & ~w16130;
assign w16159 = w11766 & w12365;
assign w16160 = ~w16157 & w16159;
assign w16161 = ~w16158 & w16160;
assign w16162 = ~w16156 & w16161;
assign w16163 = w11766 & ~w12423;
assign w16164 = w16133 & ~w16163;
assign w16165 = ~w11559 & ~w16164;
assign w16166 = ~w11635 & ~w16165;
assign w16167 = ~w16162 & w16166;
assign w16168 = ~w42 & w59;
assign w16169 = ~w90 & ~w62;
assign w16170 = ~w230 & w233;
assign w16171 = ~w259 & w262;
assign w16172 = ~w309 & ~w281;
assign w16173 = ~w355 & w371;
assign w16174 = ~w482 & w499;
assign w16175 = ~w529 & ~w531;
assign w16176 = ~w561 & ~w563;
assign w16177 = ~w592 & ~w594;
assign w16178 = ~w704 & w721;
assign w16179 = ~w781 & w786;
assign w16180 = ~w813 & w818;
assign w16181 = w824 & ~w850;
assign w16182 = ~w912 & ~w884;
assign w16183 = ~w949 & w953;
assign w16184 = ~w967 & w970;
assign w16185 = ~w995 & w998;
assign w16186 = ~w1041 & ~w1014;
assign w16187 = ~w1197 & ~w1170;
assign w16188 = ~w1339 & w1342;
assign w16189 = ~w1374 & w1377;
assign w16190 = ~w1398 & w1401;
assign w16191 = ~w1446 & ~w1431;
assign w16192 = ~w1608 & ~w1580;
assign w16193 = ~w1626 & w1629;
assign w16194 = ~w1652 & w1655;
assign w16195 = ~w1685 & w1688;
assign w16196 = ~w1709 & w1712;
assign w16197 = ~w1739 & w1742;
assign w16198 = ~w1782 & w1785;
assign w16199 = ~w1811 & w1814;
assign w16200 = ~w1841 & w1844;
assign w16201 = ~w1914 & ~w1916;
assign w16202 = ~w1978 & ~w1980;
assign w16203 = ~w2008 & ~w2010;
assign w16204 = ~w2070 & ~w2072;
assign w16205 = ~w2100 & ~w2102;
assign w16206 = ~w2131 & ~w2133;
assign w16207 = ~w2161 & ~w2163;
assign w16208 = ~w2196 & ~w2168;
assign w16209 = ~w2205 & w2223;
assign w16210 = ~w2258 & ~w2231;
assign w16211 = ~w2335 & w2338;
assign w16212 = ~w2364 & w2367;
assign w16213 = ~w2398 & ~w2388;
assign w16214 = ~w2427 & w2430;
assign w16215 = ~w2455 & w2458;
assign w16216 = ~w2494 & ~w2475;
assign w16217 = (~w1230 & ~w1670) | (~w1230 & w17428) | (~w1670 & w17428);
assign w16218 = ~w355 & w370;
assign w16219 = (w467 & ~w1670) | (w467 & w16824) | (~w1670 & w16824);
assign w16220 = (~w1420 & ~w1670) | (~w1420 & w17429) | (~w1670 & w17429);
assign w16221 = ~w2572 & ~w955;
assign w16222 = ~w2534 & w2539;
assign w16223 = ~w2383 & w2539;
assign w16224 = w2672 & ~w2671;
assign w16225 = w2700 & ~w2699;
assign w16226 = ~w3065 & w3068;
assign w16227 = ~w3092 & w3095;
assign w16228 = ~w3121 & w3124;
assign w16229 = ~w3149 & w3152;
assign w16230 = ~w3179 & w3182;
assign w16231 = ~w3207 & w3210;
assign w16232 = w2539 & w2387;
assign w16233 = ~w1758 & w3310;
assign w16234 = ~w2551 & w1199;
assign w16235 = ~w2564 & w3328;
assign w16236 = (w3331 & ~w1670) | (w3331 & w17430) | (~w1670 & w17430);
assign w16237 = (w404 & ~w2504) | (w404 & w16825) | (~w2504 & w16825);
assign w16238 = w2634 & w16826;
assign w16239 = w2634 & w16827;
assign w16240 = w2539 & w1920;
assign w16241 = ~w3306 & w17431;
assign w16242 = w2634 & w16828;
assign w16243 = ~w2561 & w2564;
assign w16244 = (~w2538 & w17432) | (~w2538 & w17433) | (w17432 & w17433);
assign w16245 = ~w2561 & ~w1417;
assign w16246 = w2634 & w16829;
assign w16247 = ~w3351 & w4700;
assign w16248 = w3351 & w3371;
assign w16249 = w3351 & w3361;
assign w16250 = ~w3306 & w16830;
assign w16251 = w4759 & w4691;
assign w16252 = ~w4810 & w4773;
assign w16253 = ~w4810 & w4751;
assign w16254 = w3352 & w3920;
assign w16255 = (w4852 & w17434) | (w4852 & w17435) | (w17434 & w17435);
assign w16256 = ~w4051 & ~w3743;
assign w16257 = ~w5476 & w5478;
assign w16258 = ~w4766 & w4692;
assign w16259 = ~w4810 & w4689;
assign w16260 = w3352 & w5513;
assign w16261 = ~w4810 & w4762;
assign w16262 = ~w4810 & w4786;
assign w16263 = (w4788 & w4759) | (w4788 & w17436) | (w4759 & w17436);
assign w16264 = ~w4766 & w4811;
assign w16265 = ~w3420 & w17437;
assign w16266 = ~w4810 & w4846;
assign w16267 = ~w5530 & w5468;
assign w16268 = ~w4672 & ~w4687;
assign w16269 = ~w5443 & w5464;
assign w16270 = ~w4813 & w1756;
assign w16271 = ~w4854 & w18485;
assign w16272 = w6126 & ~w4489;
assign w16273 = ~w5530 & w6131;
assign w16274 = ~w5443 & w6140;
assign w16275 = ~w5611 & w6142;
assign w16276 = w6144 & ~w1358;
assign w16277 = ~w5443 & w6153;
assign w16278 = ~w5530 & w5523;
assign w16279 = w6144 & ~w1043;
assign w16280 = ~w4672 & w6157;
assign w16281 = w5411 & ~w1949;
assign w16282 = ~w5611 & w6161;
assign w16283 = ~w5530 & w5599;
assign w16284 = (w5463 & ~w5428) | (w5463 & w16832) | (~w5428 & w16832);
assign w16285 = ~w4672 & w5598;
assign w16286 = ~w5533 & w5604;
assign w16287 = (w5600 & ~w5417) | (w5600 & w17841) | (~w5417 & w17841);
assign w16288 = (w5508 & ~w5428) | (w5508 & w16833) | (~w5428 & w16833);
assign w16289 = (w5506 & ~w5597) | (w5506 & w16834) | (~w5597 & w16834);
assign w16290 = ~w4672 & w5505;
assign w16291 = w6200 & w17438;
assign w16292 = (w5511 & ~w5417) | (w5511 & w17842) | (~w5417 & w17842);
assign w16293 = w6216 & w5529;
assign w16294 = (w5415 & ~w5597) | (w5415 & w16835) | (~w5597 & w16835);
assign w16295 = (w5413 & ~w5417) | (w5413 & w17843) | (~w5417 & w17843);
assign w16296 = (w5414 & ~w5428) | (w5414 & w16836) | (~w5428 & w16836);
assign w16297 = ~w5533 & w5409;
assign w16298 = (w5549 & ~w5428) | (w5549 & w16837) | (~w5428 & w16837);
assign w16299 = (w5552 & ~w5597) | (w5552 & w16838) | (~w5597 & w16838);
assign w16300 = ~w4672 & w5546;
assign w16301 = ~w5530 & w5548;
assign w16302 = ~w5533 & w5550;
assign w16303 = (w5551 & ~w5417) | (w5551 & w17844) | (~w5417 & w17844);
assign w16304 = ~w5545 & w6252;
assign w16305 = ~w4831 & w6258;
assign w16306 = ~w6266 & ~w6264;
assign w16307 = ~w5530 & w5448;
assign w16308 = (w5447 & ~w5428) | (w5447 & w16839) | (~w5428 & w16839);
assign w16309 = ~w4672 & ~w5431;
assign w16310 = (w5449 & ~w5597) | (w5449 & w16840) | (~w5597 & w16840);
assign w16311 = ~w4672 & w5485;
assign w16312 = ~w4705 & w18487;
assign w16313 = (w5493 & ~w5428) | (w5493 & w16841) | (~w5428 & w16841);
assign w16314 = ~w6296 & ~w6300;
assign w16315 = ~w5530 & w5567;
assign w16316 = ~w5533 & w5574;
assign w16317 = (w5569 & ~w5597) | (w5569 & w16842) | (~w5597 & w16842);
assign w16318 = ~w4672 & w5571;
assign w16319 = (w5573 & ~w5428) | (w5573 & w16843) | (~w5428 & w16843);
assign w16320 = ~w1104 & w6322;
assign w16321 = ~w4672 & w5430;
assign w16322 = (w5425 & ~w5523) | (w5425 & w16844) | (~w5523 & w16844);
assign w16323 = (w5427 & ~w5597) | (w5427 & w16845) | (~w5597 & w16845);
assign w16324 = w6355 & w17439;
assign w16325 = w6329 & w6380;
assign w16326 = (w6098 & ~w6147) | (w6098 & w17440) | (~w6147 & w17440);
assign w16327 = ~w6293 & w6394;
assign w16328 = ~w6261 & w6159;
assign w16329 = w6216 & w5528;
assign w16330 = ~w5481 & w5377;
assign w16331 = (w5224 & ~w6147) | (w5224 & w17441) | (~w6147 & w17441);
assign w16332 = ~w6293 & w6158;
assign w16333 = ~w6261 & w6160;
assign w16334 = w6375 & w18155;
assign w16335 = ~w6261 & w5631;
assign w16336 = ~w6293 & w5632;
assign w16337 = w6306 & w17442;
assign w16338 = w6343 & w6233;
assign w16339 = ~w6293 & ~w5461;
assign w16340 = (w3683 & ~w6147) | (w3683 & w17443) | (~w6147 & w17443);
assign w16341 = ~w6261 & w6341;
assign w16342 = w6232 & w16846;
assign w16343 = ~w6261 & w6280;
assign w16344 = (~w4519 & ~w6147) | (~w4519 & w17444) | (~w6147 & w17444);
assign w16345 = w6515 & w6522;
assign w16346 = ~w6261 & w6223;
assign w16347 = w6532 & ~w6526;
assign w16348 = (w2695 & ~w6147) | (w2695 & w17445) | (~w6147 & w17445);
assign w16349 = ~w6293 & w6199;
assign w16350 = ~w6261 & w6206;
assign w16351 = (w6204 & w6221) | (w6204 & w17446) | (w6221 & w17446);
assign w16352 = w6551 & ~w6546;
assign w16353 = w6232 & w16847;
assign w16354 = ~w6261 & w6187;
assign w16355 = w6233 & ~w6246;
assign w16356 = ~w6293 & w6239;
assign w16357 = (w2444 & ~w6147) | (w2444 & w17447) | (~w6147 & w17447);
assign w16358 = ~w6617 & ~w6616;
assign w16359 = ~w6261 & w6619;
assign w16360 = ~w6631 & w6327;
assign w16361 = w6233 & w6313;
assign w16362 = ~w6261 & w6315;
assign w16363 = ~w6293 & w6320;
assign w16364 = ~w6293 & w6130;
assign w16365 = (~w7119 & ~w6147) | (~w7119 & w17448) | (~w6147 & w17448);
assign w16366 = ~w6261 & w7139;
assign w16367 = ~w6293 & w7141;
assign w16368 = w5645 & ~w659;
assign w16369 = w6147 & w17449;
assign w16370 = (w7165 & ~w16352) | (w7165 & w17450) | (~w16352 & w17450);
assign w16371 = ~w7171 & w6382;
assign w16372 = (w6580 & ~w6438) | (w6580 & w16848) | (~w6438 & w16848);
assign w16373 = ~w6627 & w7187;
assign w16374 = (w7194 & ~w6445) | (w7194 & w17451) | (~w6445 & w17451);
assign w16375 = ~w6627 & w6406;
assign w16376 = ~w7171 & w6454;
assign w16377 = (w6448 & ~w6438) | (w6448 & w16849) | (~w6438 & w16849);
assign w16378 = ~w6627 & w7122;
assign w16379 = (w7120 & ~w6438) | (w7120 & w16850) | (~w6438 & w16850);
assign w16380 = (w7115 & ~w16352) | (w7115 & w17452) | (~w16352 & w17452);
assign w16381 = (w7119 & ~w6445) | (w7119 & w17453) | (~w6445 & w17453);
assign w16382 = (w7148 & ~w6445) | (w7148 & w17454) | (~w6445 & w17454);
assign w16383 = (~w6219 & ~w16352) | (~w6219 & w17455) | (~w16352 & w17455);
assign w16384 = ~w7171 & w7136;
assign w16385 = (w7631 & ~w6438) | (w7631 & w16851) | (~w6438 & w16851);
assign w16386 = ~w7171 & w6383;
assign w16387 = ~w6627 & w6407;
assign w16388 = ~w7171 & w6421;
assign w16389 = (w6422 & ~w16352) | (w6422 & w17456) | (~w16352 & w17456);
assign w16390 = ~w6446 & w6419;
assign w16391 = ~w6627 & w6429;
assign w16392 = w7692 & ~w7677;
assign w16393 = ~w6627 & w6502;
assign w16394 = (w6473 & ~w6438) | (w6473 & w17457) | (~w6438 & w17457);
assign w16395 = (w6476 & ~w6445) | (w6476 & w17458) | (~w6445 & w17458);
assign w16396 = (w6469 & ~w16352) | (w6469 & w17459) | (~w16352 & w17459);
assign w16397 = ~w6627 & w6489;
assign w16398 = (w6524 & ~w16352) | (w6524 & w17460) | (~w16352 & w17460);
assign w16399 = ~w6627 & w6528;
assign w16400 = ~w7171 & w6535;
assign w16401 = (w6545 & ~w6445) | (w6545 & w17461) | (~w6445 & w17461);
assign w16402 = ~w6392 & w2695;
assign w16403 = (w6611 & ~w6445) | (w6611 & w17462) | (~w6445 & w17462);
assign w16404 = ~w7171 & w6608;
assign w16405 = (w6597 & ~w6438) | (w6597 & w16852) | (~w6438 & w16852);
assign w16406 = (w6560 & ~w6445) | (w6560 & w17463) | (~w6445 & w17463);
assign w16407 = ~w7171 & w6570;
assign w16408 = ~w6627 & w6578;
assign w16409 = (w6581 & ~w6438) | (w6581 & w17464) | (~w6438 & w17464);
assign w16410 = (w6568 & ~w16352) | (w6568 & w17465) | (~w16352 & w17465);
assign w16411 = (w6639 & ~w6438) | (w6639 & w16853) | (~w6438 & w16853);
assign w16412 = (w7197 & ~w7778) | (w7197 & w16854) | (~w7778 & w16854);
assign w16413 = (w7199 & ~w7711) | (w7199 & w16855) | (~w7711 & w16855);
assign w16414 = w7881 & w17466;
assign w16415 = (w7164 & ~w7598) | (w7164 & w18090) | (~w7598 & w18090);
assign w16416 = ~w7622 & w7193;
assign w16417 = (w7219 & ~w7778) | (w7219 & w16856) | (~w7778 & w16856);
assign w16418 = (w7213 & w16857) | (w7213 & ~w7711) | (w16857 & ~w7711);
assign w16419 = (w7587 & ~w7778) | (w7587 & w16858) | (~w7778 & w16858);
assign w16420 = (w7636 & ~w7778) | (w7636 & w16859) | (~w7778 & w16859);
assign w16421 = ~w7622 & ~w7192;
assign w16422 = (w7196 & ~w7778) | (w7196 & w16860) | (~w7778 & w16860);
assign w16423 = (w8414 & ~w7711) | (w8414 & w16861) | (~w7711 & w16861);
assign w16424 = (w7650 & w16862) | (w7650 & ~w7711) | (w16862 & ~w7711);
assign w16425 = (w7683 & ~w7598) | (w7683 & w18091) | (~w7598 & w18091);
assign w16426 = (~w6523 & w16863) | (~w6523 & ~w7711) | (w16863 & ~w7711);
assign w16427 = (w7742 & ~w7778) | (w7742 & w16864) | (~w7778 & w16864);
assign w16428 = (w7737 & w16865) | (w7737 & ~w7711) | (w16865 & ~w7711);
assign w16429 = (w7716 & ~w7778) | (w7716 & w16866) | (~w7778 & w16866);
assign w16430 = (w7800 & ~w7778) | (w7800 & w16867) | (~w7778 & w16867);
assign w16431 = (w7812 & w16868) | (w7812 & ~w7711) | (w16868 & ~w7711);
assign w16432 = (w8591 & ~w7778) | (w8591 & w16869) | (~w7778 & w16869);
assign w16433 = (w7762 & ~w7598) | (w7762 & w18092) | (~w7598 & w18092);
assign w16434 = (w7777 & ~w7711) | (w7777 & w16870) | (~w7711 & w16870);
assign w16435 = ~w7622 & w7765;
assign w16436 = (w7902 & ~w7778) | (w7902 & w16871) | (~w7778 & w16871);
assign w16437 = ~w7622 & w7908;
assign w16438 = (w7910 & ~w7598) | (w7910 & w18156) | (~w7598 & w18156);
assign w16439 = (w7924 & w16872) | (w7924 & ~w7711) | (w16872 & ~w7711);
assign w16440 = (w7870 & w16873) | (w7870 & ~w7711) | (w16873 & ~w7711);
assign w16441 = (w7871 & ~w7778) | (w7871 & w16874) | (~w7778 & w16874);
assign w16442 = (w7866 & ~w7598) | (w7866 & w18093) | (~w7598 & w18093);
assign w16443 = ~w7622 & w7865;
assign w16444 = (w7846 & w16875) | (w7846 & ~w7711) | (w16875 & ~w7711);
assign w16445 = ~w7622 & w7835;
assign w16446 = (w7845 & ~w7778) | (w7845 & w16876) | (~w7778 & w16876);
assign w16447 = w8342 & ~w2011;
assign w16448 = (w8031 & w7993) | (w8031 & w17467) | (w7993 & w17467);
assign w16449 = ~w8318 & w8294;
assign w16450 = ~w6521 & w9040;
assign w16451 = ~w7585 & w7259;
assign w16452 = ~w1756 & w9047;
assign w16453 = (w8419 & ~w7987) | (w8419 & w17917) | (~w7987 & w17917);
assign w16454 = ~w1756 & w8413;
assign w16455 = ~w6521 & w8415;
assign w16456 = ~w7989 & w8367;
assign w16457 = ~w1756 & w8370;
assign w16458 = ~w6521 & w8371;
assign w16459 = ~w6521 & w7963;
assign w16460 = ~w1756 & w7961;
assign w16461 = ~w1756 & w8395;
assign w16462 = ~w6521 & w8396;
assign w16463 = w8344 & ~w5341;
assign w16464 = (w8392 & ~w7987) | (w8392 & w17918) | (~w7987 & w17918);
assign w16465 = ~w6521 & w8349;
assign w16466 = ~w1756 & w8338;
assign w16467 = w8340 & w3048;
assign w16468 = ~w1756 & w8329;
assign w16469 = ~w6521 & w8325;
assign w16470 = w8342 & ~w2164;
assign w16471 = ~w6521 & w8455;
assign w16472 = ~w1756 & w8470;
assign w16473 = (w8454 & ~w7987) | (w8454 & w17919) | (~w7987 & w17919);
assign w16474 = (w8482 & ~w7987) | (w8482 & w17920) | (~w7987 & w17920);
assign w16475 = ~w8326 & w9257;
assign w16476 = ~w1756 & w8471;
assign w16477 = ~w7989 & w8611;
assign w16478 = ~w6521 & w8604;
assign w16479 = w7979 & w3743;
assign w16480 = ~w9266 & w8514;
assign w16481 = ~w1756 & w8500;
assign w16482 = ~w8504 & ~w8499;
assign w16483 = w9317 & ~w9313;
assign w16484 = w8326 & w4313;
assign w16485 = w8340 & w2753;
assign w16486 = ~w1756 & w8518;
assign w16487 = ~w6521 & w9039;
assign w16488 = ~w7989 & w8519;
assign w16489 = ~w9327 & w18157;
assign w16490 = ~w7648 & ~w3019;
assign w16491 = w8344 & w3197;
assign w16492 = ~w7989 & w8572;
assign w16493 = ~w1756 & w8571;
assign w16494 = ~w6521 & w8693;
assign w16495 = ~w1756 & w8691;
assign w16496 = ~w7989 & w8692;
assign w16497 = w9428 & w8715;
assign w16498 = ~w1756 & w9437;
assign w16499 = w9010 & w1329;
assign w16500 = ~w6521 & w8633;
assign w16501 = w8340 & ~w1012;
assign w16502 = w7980 & w1358;
assign w16503 = w8326 & ~w1261;
assign w16504 = ~w7989 & w8635;
assign w16505 = w8344 & ~w913;
assign w16506 = ~w7989 & w8671;
assign w16507 = ~w1756 & w8670;
assign w16508 = ~w7989 & w8418;
assign w16509 = w8347 & w217;
assign w16510 = w8342 & ~w1981;
assign w16511 = w9010 & ~w5680;
assign w16512 = w8344 & ~w4895;
assign w16513 = w7648 & w9556;
assign w16514 = ~w8319 & ~w8203;
assign w16515 = ~w9433 & w9629;
assign w16516 = (w9632 & ~w9396) | (w9632 & w17468) | (~w9396 & w17468);
assign w16517 = ~w9647 & w9649;
assign w16518 = w9543 & ~w6930;
assign w16519 = (~w8051 & ~w9564) | (~w8051 & w16877) | (~w9564 & w16877);
assign w16520 = w9042 & w7317;
assign w16521 = ~w9009 & w9667;
assign w16522 = ~w9433 & w9550;
assign w16523 = (w9393 & w17469) | (w9393 & w17470) | (w17469 & w17470);
assign w16524 = w9042 & w7259;
assign w16525 = (w9030 & ~w9396) | (w9030 & w17471) | (~w9396 & w17471);
assign w16526 = (w9032 & ~w9564) | (w9032 & w18158) | (~w9564 & w18158);
assign w16527 = ~w9647 & w9024;
assign w16528 = ~w9433 & w9008;
assign w16529 = w9543 & ~w7057;
assign w16530 = ~w8319 & w8114;
assign w16531 = ~w9433 & w9095;
assign w16532 = w9222 & ~w1168;
assign w16533 = ~w9647 & w9171;
assign w16534 = ~w9647 & w9062;
assign w16535 = ~w9433 & w9061;
assign w16536 = ~w9060 & w9771;
assign w16537 = (w9213 & ~w9396) | (w9213 & w17472) | (~w9396 & w17472);
assign w16538 = ~w9433 & w9007;
assign w16539 = ~w9195 & w9069;
assign w16540 = w9817 & w16879;
assign w16541 = ~w9433 & w9191;
assign w16542 = (w9184 & ~w9396) | (w9184 & w17473) | (~w9396 & w17473);
assign w16543 = (w9185 & ~w9509) | (w9185 & w18448) | (~w9509 & w18448);
assign w16544 = ~w9647 & w9249;
assign w16545 = ~w9195 & w9253;
assign w16546 = (w9342 & ~w9564) | (w9342 & w16880) | (~w9564 & w16880);
assign w16547 = w9543 & w4342;
assign w16548 = w9060 & ~w4400;
assign w16549 = w9543 & w3595;
assign w16550 = w9441 & w3654;
assign w16551 = ~w9950 & ~w9954;
assign w16552 = ~w9195 & w9366;
assign w16553 = w9009 & ~w3019;
assign w16554 = ~w9433 & w9376;
assign w16555 = (w9991 & ~w9396) | (w9991 & w17474) | (~w9396 & w17474);
assign w16556 = ~w9195 & w9423;
assign w16557 = w9116 & w2444;
assign w16558 = (w9417 & ~w9509) | (w9417 & w18449) | (~w9509 & w18449);
assign w16559 = w10039 & w16881;
assign w16560 = ~w9565 & w9456;
assign w16561 = (w9448 & ~w9396) | (w9448 & w17475) | (~w9396 & w17475);
assign w16562 = ~w9459 & w10076;
assign w16563 = ~w9565 & w9479;
assign w16564 = (w9489 & ~w9396) | (w9489 & w17476) | (~w9396 & w17476);
assign w16565 = ~w9433 & w9486;
assign w16566 = ~w9195 & w9488;
assign w16567 = ~w9647 & w10107;
assign w16568 = ~w9647 & w9118;
assign w16569 = ~w9433 & w9121;
assign w16570 = ~w9116 & w10163;
assign w16571 = (w9123 & ~w9564) | (w9123 & w18159) | (~w9564 & w18159);
assign w16572 = (w9115 & ~w9396) | (w9115 & w17477) | (~w9396 & w17477);
assign w16573 = ~w9476 & w9167;
assign w16574 = ~w9433 & w9169;
assign w16575 = ~w9647 & w9172;
assign w16576 = ~w9027 & ~w3623;
assign w16577 = (w9149 & ~w9396) | (w9149 & w17478) | (~w9396 & w17478);
assign w16578 = w9441 & ~w5709;
assign w16579 = ~w9060 & w10262;
assign w16580 = ~w9781 & w9660;
assign w16581 = w9654 & ~w6842;
assign w16582 = ~w9963 & w10516;
assign w16583 = (w10518 & ~w10042) | (w10518 & w16882) | (~w10042 & w16882);
assign w16584 = w9627 & ~w8232;
assign w16585 = (w10522 & ~w9880) | (w10522 & w16883) | (~w9880 & w16883);
assign w16586 = (w10525 & ~w9897) | (w10525 & w18160) | (~w9897 & w18160);
assign w16587 = w10116 & w10128;
assign w16588 = ~w10007 & w10530;
assign w16589 = (w9658 & ~w10059) | (w9658 & w16884) | (~w10059 & w16884);
assign w16590 = (w10547 & ~w9823) | (w10547 & w16885) | (~w9823 & w16885);
assign w16591 = (w9634 & ~w9749) | (w9634 & w16886) | (~w9749 & w16886);
assign w16592 = ~w10544 & ~w10543;
assign w16593 = (w10201 & ~w9880) | (w10201 & w16887) | (~w9880 & w16887);
assign w16594 = (w9796 & ~w10042) | (w9796 & w16888) | (~w10042 & w16888);
assign w16595 = ~w9963 & w9900;
assign w16596 = (w9817 & ~w9823) | (w9817 & w16889) | (~w9823 & w16889);
assign w16597 = w9654 & ~w6871;
assign w16598 = (~w9363 & ~w9897) | (~w9363 & w18161) | (~w9897 & w18161);
assign w16599 = ~w10589 & w10591;
assign w16600 = (w10256 & ~w10042) | (w10256 & w16890) | (~w10042 & w16890);
assign w16601 = (w10259 & ~w9880) | (w10259 & w16891) | (~w9880 & w16891);
assign w16602 = ~w9963 & w10257;
assign w16603 = (w10260 & ~w10059) | (w10260 & w16892) | (~w10059 & w16892);
assign w16604 = (w10253 & ~w9897) | (w10253 & w18162) | (~w9897 & w18162);
assign w16605 = ~w10007 & w10254;
assign w16606 = ~w9781 & w10255;
assign w16607 = w10621 & w10555;
assign w16608 = w10202 & w9812;
assign w16609 = ~w10051 & w9984;
assign w16610 = (w9979 & ~w10225) | (w9979 & w18163) | (~w10225 & w18163);
assign w16611 = ~w10830 & w18164;
assign w16612 = w10824 & w16893;
assign w16613 = (w10019 & ~w9897) | (w10019 & w18165) | (~w9897 & w18165);
assign w16614 = (w10010 & ~w9749) | (w10010 & w18166) | (~w9749 & w18166);
assign w16615 = w9654 & w2134;
assign w16616 = ~w9963 & w10031;
assign w16617 = (~w9434 & ~w10042) | (~w9434 & w16894) | (~w10042 & w16894);
assign w16618 = (w10032 & ~w9880) | (w10032 & w18167) | (~w9880 & w18167);
assign w16619 = ~w10007 & w10018;
assign w16620 = ~w9781 & w10012;
assign w16621 = (w10011 & ~w10225) | (w10011 & w18168) | (~w10225 & w18168);
assign w16622 = ~w10868 & ~w10869;
assign w16623 = w10888 & w10898;
assign w16624 = w10126 & w18169;
assign w16625 = ~w9781 & w10124;
assign w16626 = ~w9963 & w10096;
assign w16627 = (w9701 & ~w10225) | (w9701 & w17479) | (~w10225 & w17479);
assign w16628 = ~w10099 & w10938;
assign w16629 = ~w10927 & ~w10930;
assign w16630 = w10944 & w16896;
assign w16631 = ~w9781 & w10061;
assign w16632 = w9627 & ~w1727;
assign w16633 = (w10060 & ~w9880) | (w10060 & w18170) | (~w9880 & w18170);
assign w16634 = (w9950 & ~w9823) | (w9950 & w16897) | (~w9823 & w16897);
assign w16635 = (w9955 & ~w10042) | (w9955 & w18171) | (~w10042 & w18171);
assign w16636 = (w9953 & ~w10059) | (w9953 & w18172) | (~w10059 & w18172);
assign w16637 = ~w9781 & w9936;
assign w16638 = w10128 & w18173;
assign w16639 = ~w9781 & w9886;
assign w16640 = (w9910 & ~w10225) | (w9910 & w18174) | (~w10225 & w18174);
assign w16641 = ~w9750 & w9905;
assign w16642 = (w9885 & ~w10042) | (w9885 & w18175) | (~w10042 & w18175);
assign w16643 = ~w10007 & w9888;
assign w16644 = ~w10007 & w9789;
assign w16645 = ~w9963 & w9790;
assign w16646 = ~w10552 & w16898;
assign w16647 = (w9795 & ~w10225) | (w9795 & w18176) | (~w10225 & w18176);
assign w16648 = ~w9781 & w9787;
assign w16649 = w11115 & w16899;
assign w16650 = (w9832 & ~w9880) | (w9832 & w16900) | (~w9880 & w16900);
assign w16651 = (w9827 & ~w10042) | (w9827 & w16901) | (~w10042 & w16901);
assign w16652 = ~w9963 & w9833;
assign w16653 = (w9829 & ~w10059) | (w9829 & w16902) | (~w10059 & w16902);
assign w16654 = ~w10007 & w9828;
assign w16655 = (w9830 & ~w9897) | (w9830 & w18177) | (~w9897 & w18177);
assign w16656 = (w9856 & ~w9897) | (w9856 & w18178) | (~w9897 & w18178);
assign w16657 = w9654 & w5253;
assign w16658 = (w9878 & ~w10059) | (w9878 & w18179) | (~w10059 & w18179);
assign w16659 = (w9849 & ~w10225) | (w9849 & w18180) | (~w10225 & w18180);
assign w16660 = (w9847 & ~w9749) | (w9847 & w18181) | (~w9749 & w18181);
assign w16661 = ~w9750 & w9769;
assign w16662 = w9656 & ~w7347;
assign w16663 = w9627 & ~w7259;
assign w16664 = ~w9963 & w9755;
assign w16665 = ~w10007 & w9763;
assign w16666 = (w9761 & ~w10059) | (w9761 & w16903) | (~w10059 & w16903);
assign w16667 = (w9767 & ~w9880) | (w9767 & w16904) | (~w9880 & w16904);
assign w16668 = (w9758 & ~w9897) | (w9758 & w18182) | (~w9897 & w18182);
assign w16669 = (w9762 & ~w9823) | (w9762 & w16905) | (~w9823 & w16905);
assign w16670 = ~w9781 & w11231;
assign w16671 = (w10211 & ~w10042) | (w10211 & w18183) | (~w10042 & w18183);
assign w16672 = ~w10007 & w10216;
assign w16673 = (w10213 & ~w9897) | (w10213 & w18184) | (~w9897 & w18184);
assign w16674 = (w10212 & ~w9880) | (w10212 & w18185) | (~w9880 & w18185);
assign w16675 = (w10160 & ~w10042) | (w10160 & w18186) | (~w10042 & w18186);
assign w16676 = ~w10007 & w10180;
assign w16677 = ~w9963 & w10179;
assign w16678 = (w10155 & ~w10225) | (w10155 & w18187) | (~w10225 & w18187);
assign w16679 = ~w9781 & w10156;
assign w16680 = (w10154 & ~w9749) | (w10154 & w18188) | (~w9749 & w18188);
assign w16681 = (w10158 & ~w9880) | (w10158 & w18189) | (~w9880 & w18189);
assign w16682 = (w10178 & ~w10059) | (w10178 & w18190) | (~w10059 & w18190);
assign w16683 = ~w11276 & ~w11282;
assign w16684 = w11302 & w11305;
assign w16685 = (w10202 & ~w9880) | (w10202 & w16906) | (~w9880 & w16906);
assign w16686 = (w10191 & ~w10042) | (w10191 & w16907) | (~w10042 & w16907);
assign w16687 = (w9709 & ~w9823) | (w9709 & w16908) | (~w9823 & w16908);
assign w16688 = ~w9963 & w9706;
assign w16689 = (w9708 & ~w9897) | (w9708 & w17845) | (~w9897 & w17845);
assign w16690 = (w9703 & w9968) | (w9703 & w18191) | (w9968 & w18191);
assign w16691 = (w9711 & ~w10042) | (w9711 & w16909) | (~w10042 & w16909);
assign w16692 = w9627 & w11350;
assign w16693 = ~w10007 & w9737;
assign w16694 = (w9732 & ~w9897) | (w9732 & w18192) | (~w9897 & w18192);
assign w16695 = (w9735 & ~w10042) | (w9735 & w18193) | (~w10042 & w18193);
assign w16696 = (w9736 & ~w9880) | (w9736 & w18194) | (~w9880 & w18194);
assign w16697 = (w9739 & ~w10059) | (w9739 & w18195) | (~w10059 & w18195);
assign w16698 = ~w10007 & w9676;
assign w16699 = ~w9781 & w9680;
assign w16700 = ~w10051 & w9674;
assign w16701 = ~w9881 & w9681;
assign w16702 = ~w9898 & w9673;
assign w16703 = (w9641 & ~w9823) | (w9641 & w16910) | (~w9823 & w16910);
assign w16704 = (w9650 & ~w10128) | (w9650 & w16911) | (~w10128 & w16911);
assign w16705 = (w9659 & ~w10059) | (w9659 & w16912) | (~w10059 & w16912);
assign w16706 = (w9657 & ~w9897) | (w9657 & w17846) | (~w9897 & w17846);
assign w16707 = (w9643 & ~w9962) | (w9643 & w18094) | (~w9962 & w18094);
assign w16708 = ~w10007 & w9633;
assign w16709 = (w9645 & ~w9880) | (w9645 & w16913) | (~w9880 & w16913);
assign w16710 = ~w9781 & w9661;
assign w16711 = w11432 & w10555;
assign w16712 = (w10929 & ~w11261) | (w10929 & w16914) | (~w11261 & w16914);
assign w16713 = (w10550 & ~w11406) | (w10550 & w16915) | (~w11406 & w16915);
assign w16714 = (w10551 & ~w11384) | (w10551 & w16916) | (~w11384 & w16916);
assign w16715 = (w10570 & ~w11200) | (w10570 & w16917) | (~w11200 & w16917);
assign w16716 = (w10580 & ~w11117) | (w10580 & w16918) | (~w11117 & w16918);
assign w16717 = (w10545 & ~w10964) | (w10545 & w16919) | (~w10964 & w16919);
assign w16718 = (w10572 & ~w10944) | (w10572 & w16920) | (~w10944 & w16920);
assign w16719 = (w10578 & ~w10826) | (w10578 & w16921) | (~w10826 & w16921);
assign w16720 = (w10576 & ~w11020) | (w10576 & w16922) | (~w11020 & w16922);
assign w16721 = (w10586 & ~w11067) | (w10586 & w16923) | (~w11067 & w16923);
assign w16722 = (w10512 & ~w11241) | (w10512 & w18450) | (~w11241 & w18450);
assign w16723 = (w10520 & ~w11361) | (w10520 & w18196) | (~w11361 & w18196);
assign w16724 = (w10607 & ~w11200) | (w10607 & w16924) | (~w11200 & w16924);
assign w16725 = (~w9730 & ~w11361) | (~w9730 & w18197) | (~w11361 & w18197);
assign w16726 = (~w10130 & ~w10944) | (~w10130 & w16925) | (~w10944 & w16925);
assign w16727 = (w10953 & ~w11384) | (w10953 & w16926) | (~w11384 & w16926);
assign w16728 = (w10951 & ~w10826) | (w10951 & w16927) | (~w10826 & w16927);
assign w16729 = (w10975 & ~w11020) | (w10975 & w16928) | (~w11020 & w16928);
assign w16730 = (w10976 & ~w11067) | (w10976 & w16929) | (~w11067 & w16929);
assign w16731 = (w10910 & ~w11361) | (w10910 & w18198) | (~w11361 & w18198);
assign w16732 = (w10932 & ~w11384) | (w10932 & w18199) | (~w11384 & w18199);
assign w16733 = (w10906 & ~w11241) | (w10906 & w18451) | (~w11241 & w18451);
assign w16734 = (~w9882 & ~w11200) | (~w9882 & w16930) | (~w11200 & w16930);
assign w16735 = (w10913 & ~w11117) | (w10913 & w18200) | (~w11117 & w18200);
assign w16736 = (w10911 & ~w10826) | (w10911 & w18201) | (~w10826 & w18201);
assign w16737 = (~w11066 & w18452) | (~w11066 & w18453) | (w18452 & w18453);
assign w16738 = (w10893 & ~w10944) | (w10893 & w16932) | (~w10944 & w16932);
assign w16739 = (w10866 & ~w10826) | (w10866 & w16933) | (~w10826 & w16933);
assign w16740 = (w10873 & ~w11261) | (w10873 & w16934) | (~w11261 & w16934);
assign w16741 = (w10857 & ~w11384) | (w10857 & w16935) | (~w11384 & w16935);
assign w16742 = w11829 & ~w11936;
assign w16743 = (w11031 & ~w11067) | (w11031 & w18202) | (~w11067 & w18202);
assign w16744 = (w11023 & ~w10964) | (w11023 & w18203) | (~w10964 & w18203);
assign w16745 = (w11009 & ~w11117) | (w11009 & w18204) | (~w11117 & w18204);
assign w16746 = (w11029 & ~w10826) | (w11029 & w18205) | (~w10826 & w18205);
assign w16747 = (w11028 & ~w11241) | (w11028 & w18454) | (~w11241 & w18454);
assign w16748 = (w11004 & ~w11384) | (w11004 & w16936) | (~w11384 & w16936);
assign w16749 = (w11024 & ~w11361) | (w11024 & w17847) | (~w11361 & w17847);
assign w16750 = (w11008 & ~w11261) | (w11008 & w16937) | (~w11261 & w16937);
assign w16751 = w11994 & w11993;
assign w16752 = (w7789 & ~w11020) | (w7789 & w16938) | (~w11020 & w16938);
assign w16753 = (w7786 & ~w10964) | (w7786 & w16939) | (~w10964 & w16939);
assign w16754 = (w10837 & ~w11067) | (w10837 & w16940) | (~w11067 & w16940);
assign w16755 = (w10820 & ~w10944) | (w10820 & w16941) | (~w10944 & w16941);
assign w16756 = (w10828 & ~w10964) | (w10828 & w16942) | (~w10964 & w16942);
assign w16757 = (w10835 & ~w11200) | (w10835 & w16943) | (~w11200 & w16943);
assign w16758 = (w11167 & ~w10944) | (w11167 & w16944) | (~w10944 & w16944);
assign w16759 = (w11161 & ~w11067) | (w11161 & w16945) | (~w11067 & w16945);
assign w16760 = (w11196 & ~w10826) | (w11196 & w16946) | (~w10826 & w16946);
assign w16761 = (w11197 & ~w11117) | (w11197 & w16947) | (~w11117 & w16947);
assign w16762 = (w11173 & ~w11261) | (w11173 & w16948) | (~w11261 & w16948);
assign w16763 = (w11073 & ~w10826) | (w11073 & w16949) | (~w10826 & w16949);
assign w16764 = (w11078 & ~w11200) | (w11078 & w16950) | (~w11200 & w16950);
assign w16765 = (w11052 & ~w11020) | (w11052 & w16951) | (~w11020 & w16951);
assign w16766 = (w11075 & ~w11117) | (w11075 & w16952) | (~w11117 & w16952);
assign w16767 = (w11074 & ~w10944) | (w11074 & w16953) | (~w10944 & w16953);
assign w16768 = (w11106 & ~w11406) | (w11106 & w16954) | (~w11406 & w16954);
assign w16769 = (w11129 & ~w11067) | (w11129 & w16955) | (~w11067 & w16955);
assign w16770 = (w11110 & ~w11020) | (w11110 & w16956) | (~w11020 & w16956);
assign w16771 = (w11123 & ~w11261) | (w11123 & w16957) | (~w11261 & w16957);
assign w16772 = (w11125 & ~w11241) | (w11125 & w18455) | (~w11241 & w18455);
assign w16773 = (w11128 & ~w11384) | (w11128 & w16958) | (~w11384 & w16958);
assign w16774 = (~w11066 & w18456) | (~w11066 & w18457) | (w18456 & w18457);
assign w16775 = (w11310 & ~w10964) | (w11310 & w16960) | (~w10964 & w16960);
assign w16776 = (w11313 & ~w11117) | (w11313 & w16961) | (~w11117 & w16961);
assign w16777 = (w11311 & ~w10826) | (w11311 & w16962) | (~w10826 & w16962);
assign w16778 = (w11286 & ~w11200) | (w11286 & w16963) | (~w11200 & w16963);
assign w16779 = (~w10963 & w18458) | (~w10963 & w18459) | (w18458 & w18459);
assign w16780 = (w11271 & ~w11117) | (w11271 & w16965) | (~w11117 & w16965);
assign w16781 = (w11275 & ~w10826) | (w11275 & w16966) | (~w10826 & w16966);
assign w16782 = (~w11066 & w18460) | (~w11066 & w18461) | (w18460 & w18461);
assign w16783 = (w11280 & ~w11261) | (w11280 & w16968) | (~w11261 & w16968);
assign w16784 = (w11277 & ~w11406) | (w11277 & w16969) | (~w11406 & w16969);
assign w16785 = ~w11245 & w11281;
assign w16786 = (w11278 & ~w11361) | (w11278 & w18206) | (~w11361 & w18206);
assign w16787 = ~w11245 & w11376;
assign w16788 = (w11371 & ~w11200) | (w11371 & w16970) | (~w11200 & w16970);
assign w16789 = (w11369 & ~w11020) | (w11369 & w16971) | (~w11020 & w16971);
assign w16790 = (w11374 & ~w11117) | (w11374 & w16972) | (~w11117 & w16972);
assign w16791 = (w11339 & ~w11067) | (w11339 & w16973) | (~w11067 & w16973);
assign w16792 = (w11345 & ~w10964) | (w11345 & w16974) | (~w10964 & w16974);
assign w16793 = (w11344 & ~w11200) | (w11344 & w16975) | (~w11200 & w16975);
assign w16794 = (w11340 & ~w10826) | (w11340 & w16976) | (~w10826 & w16976);
assign w16795 = (w11336 & ~w11020) | (w11336 & w16977) | (~w11020 & w16977);
assign w16796 = (w11337 & ~w10944) | (w11337 & w16978) | (~w10944 & w16978);
assign w16797 = (w11335 & ~w11406) | (w11335 & w16979) | (~w11406 & w16979);
assign w16798 = (w11417 & ~w11020) | (w11417 & w16980) | (~w11020 & w16980);
assign w16799 = (w11415 & ~w11067) | (w11415 & w16981) | (~w11067 & w16981);
assign w16800 = (w11414 & ~w10964) | (w11414 & w16982) | (~w10964 & w16982);
assign w16801 = (w11412 & ~w11117) | (w11412 & w16983) | (~w11117 & w16983);
assign w16802 = (w11419 & ~w11200) | (w11419 & w16984) | (~w11200 & w16984);
assign w16803 = (w11418 & ~w10826) | (w11418 & w16985) | (~w10826 & w16985);
assign w16804 = (w11413 & ~w10944) | (w11413 & w16986) | (~w10944 & w16986);
assign w16805 = (w11397 & ~w10964) | (w11397 & w16987) | (~w10964 & w16987);
assign w16806 = (w11395 & ~w11067) | (w11395 & w16988) | (~w11067 & w16988);
assign w16807 = (w11394 & ~w11200) | (w11394 & w16989) | (~w11200 & w16989);
assign w16808 = (w11399 & ~w11117) | (w11399 & w16990) | (~w11117 & w16990);
assign w16809 = (w11390 & ~w11361) | (w11390 & w18207) | (~w11361 & w18207);
assign w16810 = (w11389 & ~w10826) | (w11389 & w18208) | (~w10826 & w18208);
assign w16811 = (w11223 & ~w11067) | (w11223 & w18209) | (~w11067 & w18209);
assign w16812 = (w11221 & ~w10964) | (w11221 & w18210) | (~w10964 & w18210);
assign w16813 = (w11212 & ~w11384) | (w11212 & w18211) | (~w11384 & w18211);
assign w16814 = (w11226 & ~w11117) | (w11226 & w18212) | (~w11117 & w18212);
assign w16815 = (w11219 & ~w11020) | (w11219 & w18213) | (~w11020 & w18213);
assign w16816 = (w11220 & ~w10826) | (w11220 & w18214) | (~w10826 & w18214);
assign w16817 = ~w11042 & w11256;
assign w16818 = w12330 & pi022;
assign w16819 = w12327 & pi020;
assign w16820 = w11480 & pi023;
assign w16821 = w12330 & pi021;
assign w16822 = ~w16141 & w16131;
assign w16823 = w15523 & ~w11996;
assign w16824 = ~w1756 & w467;
assign w16825 = ~w2535 & w404;
assign w16826 = ~w342 & ~w1012;
assign w16827 = ~w342 & w2383;
assign w16828 = ~w342 & w3054;
assign w16829 = ~w342 & ~w3258;
assign w16830 = w2586 & ~w373;
assign w16831 = ~w4744 & w5424;
assign w16832 = ~w16255 & w5463;
assign w16833 = ~w16255 & w5508;
assign w16834 = ~w4839 & w5506;
assign w16835 = ~w4839 & w5415;
assign w16836 = ~w16255 & w5414;
assign w16837 = ~w16255 & w5549;
assign w16838 = ~w4839 & w5552;
assign w16839 = ~w16255 & w5447;
assign w16840 = ~w4839 & w5449;
assign w16841 = ~w16255 & w5493;
assign w16842 = ~w4839 & w5569;
assign w16843 = ~w16255 & w5573;
assign w16844 = ~w5529 & w5425;
assign w16845 = ~w4839 & w5427;
assign w16846 = ~w3287 & w6222;
assign w16847 = ~w3287 & w6186;
assign w16848 = w6427 & w6580;
assign w16849 = w6427 & w6448;
assign w16850 = w6427 & w7120;
assign w16851 = w6427 & w7631;
assign w16852 = w6427 & w6597;
assign w16853 = w6427 & w6639;
assign w16854 = ~w7781 & w7197;
assign w16855 = ~w7752 & w7199;
assign w16856 = ~w7781 & w7219;
assign w16857 = ~w7752 & w7213;
assign w16858 = ~w7781 & w7587;
assign w16859 = ~w7781 & w7636;
assign w16860 = ~w7781 & w7196;
assign w16861 = ~w7752 & w8414;
assign w16862 = ~w7752 & w7650;
assign w16863 = ~w7752 & ~w6523;
assign w16864 = ~w7781 & w7742;
assign w16865 = ~w7752 & w7737;
assign w16866 = ~w7781 & w7716;
assign w16867 = ~w7781 & w7800;
assign w16868 = ~w7752 & w7812;
assign w16869 = ~w7781 & w8591;
assign w16870 = ~w7752 & w7777;
assign w16871 = ~w7781 & w7902;
assign w16872 = ~w7752 & w7924;
assign w16873 = ~w7752 & w7870;
assign w16874 = ~w7781 & w7871;
assign w16875 = ~w7752 & w7846;
assign w16876 = ~w7781 & w7845;
assign w16877 = w9555 & ~w8051;
assign w16878 = ~w7806 & w9183;
assign w16879 = w6037 & w5949;
assign w16880 = w9555 & w9342;
assign w16881 = (w10050 & w9058) | (w10050 & w18215) | (w9058 & w18215);
assign w16882 = ~w16559 & w10518;
assign w16883 = ~w8462 & w10522;
assign w16884 = ~w9438 & w9658;
assign w16885 = ~w16540 & w10547;
assign w16886 = (w17267 & w18216) | (w17267 & w18217) | (w18216 & w18217);
assign w16887 = ~w8462 & w10201;
assign w16888 = ~w16559 & w9796;
assign w16889 = ~w16540 & w9817;
assign w16890 = ~w16559 & w10256;
assign w16891 = ~w8462 & w10259;
assign w16892 = ~w9438 & w10260;
assign w16893 = (w9971 & w10527) | (w9971 & w10007) | (w10527 & w10007);
assign w16894 = (~w9434 & ~w10039) | (~w9434 & w18218) | (~w10039 & w18218);
assign w16895 = w9171 & w10902;
assign w16896 = w7892 & w10947;
assign w16897 = ~w16540 & w9950;
assign w16898 = ~w8499 & ~w9816;
assign w16899 = (~w5889 & w10527) | (~w5889 & w18219) | (w10527 & w18219);
assign w16900 = ~w8462 & w9832;
assign w16901 = ~w16559 & w9827;
assign w16902 = ~w9438 & w9829;
assign w16903 = ~w9438 & w9761;
assign w16904 = ~w8462 & w9767;
assign w16905 = ~w16540 & w9762;
assign w16906 = ~w8462 & w10202;
assign w16907 = ~w16559 & w10191;
assign w16908 = ~w16540 & w9709;
assign w16909 = (w9711 & ~w10039) | (w9711 & w18220) | (~w10039 & w18220);
assign w16910 = ~w16540 & w9641;
assign w16911 = ~w9171 & w9650;
assign w16912 = ~w9438 & w9659;
assign w16913 = ~w8462 & w9645;
assign w16914 = w11256 & w10929;
assign w16915 = w11399 & w10550;
assign w16916 = w11374 & w10551;
assign w16917 = ~w11201 & w10570;
assign w16918 = (w10580 & ~w11115) | (w10580 & w18221) | (~w11115 & w18221);
assign w16919 = ~w10988 & w10545;
assign w16920 = ~w9015 & w10572;
assign w16921 = (w10578 & ~w10824) | (w10578 & w18222) | (~w10824 & w18222);
assign w16922 = ~w9931 & w10576;
assign w16923 = ~w9899 & w10586;
assign w16924 = ~w11201 & w10607;
assign w16925 = ~w9015 & ~w10130;
assign w16926 = w11374 & w10953;
assign w16927 = (w10951 & ~w10824) | (w10951 & w18223) | (~w10824 & w18223);
assign w16928 = ~w9931 & w10975;
assign w16929 = ~w9899 & w10976;
assign w16930 = ~w11201 & ~w9882;
assign w16931 = ~w9899 & w10856;
assign w16932 = ~w9015 & w10893;
assign w16933 = (w10866 & ~w10824) | (w10866 & w18224) | (~w10824 & w18224);
assign w16934 = w11256 & w10873;
assign w16935 = w10580 & w18225;
assign w16936 = w11374 & w11004;
assign w16937 = w11256 & w11008;
assign w16938 = ~w9931 & w7789;
assign w16939 = ~w10988 & w7786;
assign w16940 = ~w9899 & w10837;
assign w16941 = ~w9015 & w10820;
assign w16942 = ~w10988 & w10828;
assign w16943 = ~w11201 & w10835;
assign w16944 = ~w9015 & w11167;
assign w16945 = ~w9899 & w11161;
assign w16946 = (w11196 & ~w10824) | (w11196 & w18226) | (~w10824 & w18226);
assign w16947 = ~w16649 & w11197;
assign w16948 = w11256 & w11173;
assign w16949 = ~w16612 & w11073;
assign w16950 = ~w11201 & w11078;
assign w16951 = ~w9931 & w11052;
assign w16952 = ~w16649 & w11075;
assign w16953 = ~w9015 & w11074;
assign w16954 = w11399 & w11106;
assign w16955 = ~w9899 & w11129;
assign w16956 = ~w9931 & w11110;
assign w16957 = w11256 & w11123;
assign w16958 = w11374 & w11128;
assign w16959 = ~w9899 & w11151;
assign w16960 = ~w10988 & w11310;
assign w16961 = ~w16649 & w11313;
assign w16962 = ~w16612 & w11311;
assign w16963 = ~w11201 & w11286;
assign w16964 = ~w10988 & w11287;
assign w16965 = (w11271 & ~w11115) | (w11271 & w18227) | (~w11115 & w18227);
assign w16966 = (w11275 & ~w10824) | (w11275 & w18228) | (~w10824 & w18228);
assign w16967 = ~w9899 & w11276;
assign w16968 = w11256 & w11280;
assign w16969 = w11399 & w11277;
assign w16970 = ~w11201 & w11371;
assign w16971 = ~w9931 & w11369;
assign w16972 = ~w16649 & w11374;
assign w16973 = ~w9899 & w11339;
assign w16974 = ~w10988 & w11345;
assign w16975 = ~w11201 & w11344;
assign w16976 = (w11340 & ~w10824) | (w11340 & w18229) | (~w10824 & w18229);
assign w16977 = ~w9931 & w11336;
assign w16978 = ~w9015 & w11337;
assign w16979 = w11399 & w11335;
assign w16980 = ~w9931 & w11417;
assign w16981 = ~w9899 & w11415;
assign w16982 = ~w10988 & w11414;
assign w16983 = (w11412 & ~w11115) | (w11412 & w18230) | (~w11115 & w18230);
assign w16984 = ~w11201 & w11419;
assign w16985 = (w11418 & ~w10824) | (w11418 & w18231) | (~w10824 & w18231);
assign w16986 = ~w9015 & w11413;
assign w16987 = ~w10988 & w11397;
assign w16988 = ~w9899 & w11395;
assign w16989 = ~w11201 & w11394;
assign w16990 = ~w16649 & w11399;
assign w16991 = ~w1450 & ~w1424;
assign w16992 = ~w1481 & ~w1453;
assign w16993 = ~w1491 & ~w1514;
assign w16994 = ~w1544 & ~w1516;
assign w16995 = ~w1633 & w1638;
assign w16996 = ~w1659 & w1662;
assign w16997 = ~w1692 & w1697;
assign w16998 = ~w1716 & w1721;
assign w16999 = ~w1746 & w1749;
assign w17000 = ~w2561 & ~w2582;
assign w17001 = ~w2587 & ~w3346;
assign w17002 = w2634 & w373;
assign w17003 = w2586 & w3313;
assign w17004 = ~w3308 & w3365;
assign w17005 = w2634 & ~w404;
assign w17006 = w2582 & ~w852;
assign w17007 = ~w4039 & w4048;
assign w17008 = ~w4049 & ~w4009;
assign w17009 = ~w3401 & w4673;
assign w17010 = ~w3405 & w4675;
assign w17011 = w4073 & ~w2632;
assign w17012 = ~w3405 & w3389;
assign w17013 = ~w3405 & w4043;
assign w17014 = ~w3401 & w4749;
assign w17015 = w4677 & ~w2260;
assign w17016 = ~w4049 & ~w4038;
assign w17017 = ~w3401 & ~w3296;
assign w17018 = ~w3405 & w4776;
assign w17019 = ~w3401 & w3372;
assign w17020 = w4073 & w3380;
assign w17021 = ~w3405 & w3373;
assign w17022 = w2502 & ~w4049;
assign w17023 = ~w4049 & w1417;
assign w17024 = ~w4821 & ~w4820;
assign w17025 = w4804 & w1950;
assign w17026 = ~w4049 & w278;
assign w17027 = w4073 & w3409;
assign w17028 = ~w3401 & w3408;
assign w17029 = ~w4833 & w17481;
assign w17030 = (~w4071 & w4770) | (~w4071 & w17848) | (w4770 & w17848);
assign w17031 = w4103 & w17482;
assign w17032 = ~w4830 & w4752;
assign w17033 = (w4745 & w4770) | (w4745 & w17849) | (w4770 & w17849);
assign w17034 = ~w4810 & w4104;
assign w17035 = ~w4756 & w4105;
assign w17036 = (w4676 & w4832) | (w4676 & w17922) | (w4832 & w17922);
assign w17037 = ~w4830 & w4679;
assign w17038 = w4103 & w17483;
assign w17039 = ~w4830 & w5465;
assign w17040 = ~w4810 & w5471;
assign w17041 = w4103 & w17484;
assign w17042 = ~w4853 & w5483;
assign w17043 = w4103 & w17485;
assign w17044 = ~w4830 & w5486;
assign w17045 = ~w4782 & ~w5488;
assign w17046 = ~w4810 & w5490;
assign w17047 = ~w4756 & w5492;
assign w17048 = w4103 & w17486;
assign w17049 = (w4696 & w4832) | (w4696 & w17487) | (w4832 & w17487);
assign w17050 = (w4695 & ~w4748) | (w4695 & w17488) | (~w4748 & w17488);
assign w17051 = ~w4830 & w4690;
assign w17052 = (w4698 & w4770) | (w4698 & w17850) | (w4770 & w17850);
assign w17053 = w4774 & ~w3197;
assign w17054 = ~w4853 & w4759;
assign w17055 = ~w4830 & w4761;
assign w17056 = w4104 & w2473;
assign w17057 = (w4793 & ~w4748) | (w4793 & w17489) | (~w4748 & w17489);
assign w17058 = (w4794 & w4770) | (w4794 & w17851) | (w4770 & w17851);
assign w17059 = (w4789 & w4832) | (w4789 & w17490) | (w4832 & w17490);
assign w17060 = ~w4853 & w5568;
assign w17061 = ~w4684 & w1292;
assign w17062 = ~w4756 & w4812;
assign w17063 = ~w4782 & w4814;
assign w17064 = w4809 & w5576;
assign w17065 = ~w4853 & w16265;
assign w17066 = w4104 & ~w754;
assign w17067 = ~w4782 & w4834;
assign w17068 = (w4833 & ~w4748) | (w4833 & w17491) | (~w4748 & w17491);
assign w17069 = w5608 & w5611;
assign w17070 = (~w5629 & ~w5474) | (~w5629 & w17852) | (~w5474 & w17852);
assign w17071 = ~w5555 & w5466;
assign w17072 = ~w5501 & ~w4742;
assign w17073 = w5474 & w17923;
assign w17074 = ~w5555 & w6133;
assign w17075 = w5474 & w17853;
assign w17076 = ~w5555 & w16281;
assign w17077 = ~w5407 & w18488;
assign w17078 = (w5474 & w17077) | (w5474 & w17924) | (w17077 & w17924);
assign w17079 = (w883 & ~w5474) | (w883 & w17854) | (~w5474 & w17854);
assign w17080 = ~w5501 & w5593;
assign w17081 = ~w5555 & w5603;
assign w17082 = (w5506 & ~w5597) | (w5506 & w17855) | (~w5597 & w17855);
assign w17083 = (w5506 & w16289) | (w5506 & ~w5608) | (w16289 & ~w5608);
assign w17084 = w16290 | w5505;
assign w17085 = (w5505 & w16290) | (w5505 & ~w5459) | (w16290 & ~w5459);
assign w17086 = ~w5501 & w5509;
assign w17087 = (~w3048 & ~w5474) | (~w3048 & w17856) | (~w5474 & w17856);
assign w17088 = ~w5555 & w5510;
assign w17089 = ~w5555 & w5412;
assign w17090 = (w5552 & ~w5597) | (w5552 & w17857) | (~w5597 & w17857);
assign w17091 = (w5552 & w16299) | (w5552 & ~w5608) | (w16299 & ~w5608);
assign w17092 = w16300 | w5546;
assign w17093 = (w5546 & w16300) | (w5546 & ~w5459) | (w16300 & ~w5459);
assign w17094 = (w2291 & ~w5474) | (w2291 & w17858) | (~w5474 & w17858);
assign w17095 = ~w5501 & w5556;
assign w17096 = ~w5555 & w16305;
assign w17097 = ~w311 & w5644;
assign w17098 = ~w311 & w16271;
assign w17099 = ~w5555 & w5536;
assign w17100 = ~w5501 & w5451;
assign w17101 = (w4163 & ~w5474) | (w4163 & w18232) | (~w5474 & w18232);
assign w17102 = ~w5555 & w5450;
assign w17103 = w16309 | ~w5431;
assign w17104 = (~w5431 & w16309) | (~w5431 & ~w5459) | (w16309 & ~w5459);
assign w17105 = (w5449 & ~w5597) | (w5449 & w18095) | (~w5597 & w18095);
assign w17106 = (w5449 & w16310) | (w5449 & ~w5608) | (w16310 & ~w5608);
assign w17107 = w16311 | w5485;
assign w17108 = (w5485 & w16311) | (w5485 & ~w5459) | (w16311 & ~w5459);
assign w17109 = ~w5555 & w5487;
assign w17110 = w6305 & w5638;
assign w17111 = ~w5501 & w5572;
assign w17112 = ~w5555 & w5566;
assign w17113 = ~w4808 & ~w5574;
assign w17114 = (~w4808 & w5533) | (~w4808 & w17113) | (w5533 & w17113);
assign w17115 = w16317 | w5569;
assign w17116 = (w5569 & w16317) | (w5569 & ~w5608) | (w16317 & ~w5608);
assign w17117 = w16318 | w5571;
assign w17118 = (w5571 & w16318) | (w5571 & ~w5459) | (w16318 & ~w5459);
assign w17119 = ~w5480 & w3743;
assign w17120 = ~w5555 & w5433;
assign w17121 = ~w5501 & w5435;
assign w17122 = w16321 | w5430;
assign w17123 = (w5430 & w16321) | (w5430 & ~w5459) | (w16321 & ~w5459);
assign w17124 = w6389 & ~w6140;
assign w17125 = w5441 & w17925;
assign w17126 = (w6398 & ~w6177) | (w6398 & w18096) | (~w6177 & w18096);
assign w17127 = (~w5481 & ~w5635) | (~w5481 & w17859) | (~w5635 & w17859);
assign w17128 = (w6162 & ~w6177) | (w6162 & w17492) | (~w6177 & w17492);
assign w17129 = w6375 & w18489;
assign w17130 = (w6443 & w16334) | (w6443 & w5636) | (w16334 & w5636);
assign w17131 = ~w6293 & w5633;
assign w17132 = (w5646 & ~w6177) | (w5646 & w18097) | (~w6177 & w18097);
assign w17133 = ~w6454 & ~w6455;
assign w17134 = w5430 & ~w5461;
assign w17135 = ~w6293 & w17134;
assign w17136 = (w6346 & ~w6177) | (w6346 & w17926) | (~w6177 & w17926);
assign w17137 = (w5424 & ~w6412) | (w5424 & w17493) | (~w6412 & w17493);
assign w17138 = w16342 | w6222;
assign w17139 = (w6222 & w16342) | (w6222 & ~w6230) | (w16342 & ~w6230);
assign w17140 = (w6279 & ~w5635) | (w6279 & w17860) | (~w5635 & w17860);
assign w17141 = w6519 & w5632;
assign w17142 = ~w6293 & w17141;
assign w17143 = (w6221 & ~w6177) | (w6221 & w17494) | (~w6177 & w17494);
assign w17144 = (w6205 & ~w5635) | (w6205 & w17927) | (~w5635 & w17927);
assign w17145 = (w6198 & ~w6177) | (w6198 & w17928) | (~w6177 & w17928);
assign w17146 = w16353 | w6186;
assign w17147 = (w6186 & w16353) | (w6186 & ~w6230) | (w16353 & ~w6230);
assign w17148 = ~w6305 & w6184;
assign w17149 = w6574 & ~w6570;
assign w17150 = (w6243 & ~w5635) | (w6243 & w17861) | (~w5635 & w17861);
assign w17151 = (w6237 & ~w6177) | (w6237 & w17495) | (~w6177 & w17495);
assign w17152 = ~w6631 & w18490;
assign w17153 = (w6634 & w16360) | (w6634 & w6178) | (w16360 & w6178);
assign w17154 = (w6311 & ~w5635) | (w6311 & w17862) | (~w5635 & w17862);
assign w17155 = (w6303 & ~w6177) | (w6303 & w17496) | (~w6177 & w17496);
assign w17156 = (w6143 & ~w6177) | (w6143 & w17497) | (~w6177 & w17497);
assign w17157 = (w16368 & ~w6177) | (w16368 & w18098) | (~w6177 & w18098);
assign w17158 = ~w7147 & ~w7135;
assign w17159 = (w7146 & ~w17149) | (w7146 & w17929) | (~w17149 & w17929);
assign w17160 = (~w6307 & ~w6680) | (~w6307 & w17863) | (~w6680 & w17863);
assign w17161 = ~w6493 & w7117;
assign w17162 = ~w6516 & w6450;
assign w17163 = ~w6516 & w6451;
assign w17164 = (w6412 & ~w17133) | (w6412 & w17864) | (~w17133 & w17864);
assign w17165 = (w6452 & ~w6491) | (w6452 & w17930) | (~w6491 & w17930);
assign w17166 = ~w6516 & w7142;
assign w17167 = (w7138 & ~w6491) | (w7138 & w17931) | (~w6491 & w17931);
assign w17168 = (w7147 & ~w17149) | (w7147 & w17865) | (~w17149 & w17865);
assign w17169 = ~w6493 & w7635;
assign w17170 = w3019 & w7165;
assign w17171 = (w3019 & ~w6542) | (w3019 & w17498) | (~w6542 & w17498);
assign w17172 = w7152 & ~w7630;
assign w17173 = ~w6516 & w6395;
assign w17174 = (w6423 & ~w17133) | (w6423 & w17932) | (~w17133 & w17932);
assign w17175 = (w6500 & ~w6530) | (w6500 & w17499) | (~w6530 & w17499);
assign w17176 = ~w6516 & w6676;
assign w17177 = ~w2990 & w7165;
assign w17178 = (~w2990 & ~w6542) | (~w2990 & w17500) | (~w6542 & w17500);
assign w17179 = (w6673 & ~w17149) | (w6673 & w17866) | (~w17149 & w17866);
assign w17180 = (w6678 & ~w6491) | (w6678 & w17933) | (~w6491 & w17933);
assign w17181 = ~w6493 & w6527;
assign w17182 = w7793 & ~w7785;
assign w17183 = (w6544 & ~w6530) | (w6544 & w17934) | (~w6530 & w17934);
assign w17184 = ~w6516 & w6537;
assign w17185 = (w6601 & ~w6680) | (w6601 & w17935) | (~w6680 & w17935);
assign w17186 = w6241 & ~w6219;
assign w17187 = (w6241 & ~w6542) | (w6241 & w17501) | (~w6542 & w17501);
assign w17188 = ~w6493 & w6594;
assign w17189 = ~w6516 & w6598;
assign w17190 = ~w6516 & w6577;
assign w17191 = (w6569 & ~w6491) | (w6569 & w18233) | (~w6491 & w18233);
assign w17192 = (w6567 & ~w6530) | (w6567 & w17936) | (~w6530 & w17936);
assign w17193 = w7832 & w7897;
assign w17194 = (w6637 & ~w6491) | (w6637 & w18234) | (~w6491 & w18234);
assign w17195 = (w6632 & ~w17149) | (w6632 & w17937) | (~w17149 & w17937);
assign w17196 = (w6643 & ~w17133) | (w6643 & w18235) | (~w17133 & w18235);
assign w17197 = (w6640 & ~w6530) | (w6640 & w17502) | (~w6530 & w17502);
assign w17198 = ~w6516 & w6642;
assign w17199 = (w7185 & ~w7879) | (w7185 & w17867) | (~w7879 & w17867);
assign w17200 = (w7176 & ~w7693) | (w7176 & w17503) | (~w7693 & w17503);
assign w17201 = ~w7823 & w7167;
assign w17202 = (w7168 & ~w7205) | (w7168 & w17504) | (~w7205 & w17504);
assign w17203 = ~w7884 & w7215;
assign w17204 = ~w7823 & w7220;
assign w17205 = (w7225 & ~w7693) | (w7225 & w17505) | (~w7693 & w17505);
assign w17206 = ~w7823 & w7166;
assign w17207 = (w7175 & ~w7693) | (w7175 & w17506) | (~w7693 & w17506);
assign w17208 = (w7632 & ~w7693) | (w7632 & w17507) | (~w7693 & w17507);
assign w17209 = ~w7823 & w7638;
assign w17210 = ~w7694 & w7611;
assign w17211 = (w7613 & ~w7879) | (w7613 & w17868) | (~w7879 & w17868);
assign w17212 = (w8410 & ~w7879) | (w8410 & w17869) | (~w7879 & w17869);
assign w17213 = (~w7113 & ~w7205) | (~w7113 & w17508) | (~w7205 & w17508);
assign w17214 = ~w7823 & w7654;
assign w17215 = w6098 & w7164;
assign w17216 = (w6098 & ~w7599) | (w6098 & w17870) | (~w7599 & w17870);
assign w17217 = (w7651 & ~w7693) | (w7651 & w17509) | (~w7693 & w17509);
assign w17218 = (w7652 & ~w7879) | (w7652 & w17871) | (~w7879 & w17871);
assign w17219 = (w7655 & ~w7205) | (w7655 & w17510) | (~w7205 & w17510);
assign w17220 = ~w7823 & w7676;
assign w17221 = ~w7884 & w7741;
assign w17222 = ~w7823 & w7738;
assign w17223 = ~w7823 & w8563;
assign w17224 = (w7805 & ~w7879) | (w7805 & w17872) | (~w7879 & w17872);
assign w17225 = (w7813 & ~w7205) | (w7813 & w17511) | (~w7205 & w17511);
assign w17226 = w2695 & w7164;
assign w17227 = (w2695 & ~w7599) | (w2695 & w17873) | (~w7599 & w17873);
assign w17228 = (w7808 & ~w7693) | (w7808 & w17512) | (~w7693 & w17512);
assign w17229 = (w7756 & ~w7693) | (w7756 & w17513) | (~w7693 & w17513);
assign w17230 = w8599 & ~w7762;
assign w17231 = w7599 & w17874;
assign w17232 = (w7776 & ~w7879) | (w7776 & w17875) | (~w7879 & w17875);
assign w17233 = ~w7884 & w8663;
assign w17234 = (w7868 & ~w7693) | (w7868 & w17514) | (~w7693 & w17514);
assign w17235 = (w7869 & ~w7822) | (w7869 & w17876) | (~w7822 & w17876);
assign w17236 = ~w8679 & ~w8682;
assign w17237 = (w7847 & ~w7879) | (w7847 & w17877) | (~w7879 & w17877);
assign w17238 = (w7829 & ~w7205) | (w7829 & w17515) | (~w7205 & w17515);
assign w17239 = w2444 & w7164;
assign w17240 = (w2444 & ~w7599) | (w2444 & w17878) | (~w7599 & w17878);
assign w17241 = (w7841 & ~w7693) | (w7841 & w17516) | (~w7693 & w17516);
assign w17242 = w7988 & w9034;
assign w17243 = (w9044 & ~w8469) | (w9044 & w17517) | (~w8469 & w17517);
assign w17244 = (w8368 & ~w8399) | (w8368 & w18099) | (~w8399 & w18099);
assign w17245 = (w8417 & ~w8469) | (w8417 & w17518) | (~w8469 & w17518);
assign w17246 = (w8360 & ~w8469) | (w8360 & w17519) | (~w8469 & w17519);
assign w17247 = (w7983 & ~w8399) | (w7983 & w18100) | (~w8399 & w18100);
assign w17248 = (w7980 & ~w8355) | (w7980 & w17520) | (~w8355 & w17520);
assign w17249 = (w7970 & ~w8469) | (w7970 & w17521) | (~w8469 & w17521);
assign w17250 = (w8345 & ~w8469) | (w8345 & w17522) | (~w8469 & w17522);
assign w17251 = (w8440 & ~w8355) | (w8440 & w17523) | (~w8355 & w17523);
assign w17252 = (w8441 & ~w8469) | (w8441 & w17524) | (~w8469 & w17524);
assign w17253 = (w8472 & ~w8355) | (w8472 & w17525) | (~w8355 & w17525);
assign w17254 = (w8597 & ~w8469) | (w8597 & w17526) | (~w8469 & w17526);
assign w17255 = ~w8385 & ~w8391;
assign w17256 = (w8594 & ~w8355) | (w8594 & w17527) | (~w8355 & w17527);
assign w17257 = (w8526 & ~w8469) | (w8526 & w17528) | (~w8469 & w17528);
assign w17258 = (w8517 & ~w8355) | (w8517 & w17529) | (~w8355 & w17529);
assign w17259 = (w8573 & ~w8355) | (w8573 & w17530) | (~w8355 & w17530);
assign w17260 = (w8634 & ~w8469) | (w8634 & w17531) | (~w8469 & w17531);
assign w17261 = (w8680 & ~w8355) | (w8680 & w17532) | (~w8355 & w17532);
assign w17262 = (w8681 & ~w8399) | (w8681 & w18236) | (~w8399 & w18236);
assign w17263 = ~w6521 & w8667;
assign w17264 = ~w7028 & ~w7977;
assign w17265 = ~w8515 & w16512;
assign w17266 = w7626 & w9171;
assign w17267 = w7626 & ~w9504;
assign w17268 = ~w9565 & w9071;
assign w17269 = ~w9323 & w9190;
assign w17270 = ~w9433 & w9329;
assign w17271 = w9222 & ~w1292;
assign w17272 = w4163 & w9069;
assign w17273 = ~w9195 & w17272;
assign w17274 = ~w9433 & w9301;
assign w17275 = (~w9421 & w9195) | (~w9421 & w9427) | (w9195 & w9427);
assign w17276 = ~w9195 & w9455;
assign w17277 = w7903 & ~w9504;
assign w17278 = w9543 & ~w628;
assign w17279 = ~w8516 & w8384;
assign w17280 = w9543 & ~w6901;
assign w17281 = ~w8319 & w8291;
assign w17282 = w9042 & w7288;
assign w17283 = ~w9027 & ~w3449;
assign w17284 = w9547 & w91;
assign w17285 = w9146 & ~w5042;
assign w17286 = w9222 & w1699;
assign w17287 = ~w1610 & w9658;
assign w17288 = ~w1610 & w16589;
assign w17289 = ~w10272 & ~w9621;
assign w17290 = ~w10552 & w18237;
assign w17291 = w10553 & ~w16591;
assign w17292 = w9682 & w154;
assign w17293 = ~w10007 & w9675;
assign w17294 = w9627 & w8261;
assign w17295 = ~w9825 & w10246;
assign w17296 = ~w9682 & w10810;
assign w17297 = ~w1230 & w9658;
assign w17298 = ~w1230 & w16589;
assign w17299 = w2164 & w9817;
assign w17300 = w2164 & w16596;
assign w17301 = w9740 & w7847;
assign w17302 = (w10897 & w10527) | (w10897 & w18238) | (w10527 & w18238);
assign w17303 = w10989 & pi003;
assign w17304 = ~w10994 & w10996;
assign w17305 = ~w11077 & ~w11079;
assign w17306 = ~w9963 & w9319;
assign w17307 = ~w9320 & w9317;
assign w17308 = w11100 & w10552;
assign w17309 = w9816 & w10553;
assign w17310 = w10553 & ~w9812;
assign w17311 = w10553 & ~w16608;
assign w17312 = ~w5799 & w9817;
assign w17313 = ~w5799 & w16596;
assign w17314 = (w9810 & w18239) | (w9810 & w18240) | (w18239 & w18240);
assign w17315 = (w10190 & ~w10059) | (w10190 & w18241) | (~w10059 & w18241);
assign w17316 = ~w10007 & w10187;
assign w17317 = ~w10272 & w9699;
assign w17318 = ~w10272 & w9635;
assign w17319 = ~w10051 & w9630;
assign w17320 = (w10552 & ~w11099) | (w10552 & w18242) | (~w11099 & w18242);
assign w17321 = w10574 & ~w1886;
assign w17322 = w10514 & ~w6753;
assign w17323 = ~w1515 & w10545;
assign w17324 = ~w1515 & w16717;
assign w17325 = w501 & w10572;
assign w17326 = w501 & w16718;
assign w17327 = ~w2842 & w10578;
assign w17328 = ~w2842 & w16719;
assign w17329 = ~w10601 & ~w10542;
assign w17330 = ~w9672 & w9637;
assign w17331 = ~w7495 & w11516;
assign w17332 = w11520 & ~w11508;
assign w17333 = ~w9672 & w11542;
assign w17334 = w8143 & ~w11511;
assign w17335 = ~w11552 & pi027;
assign w17336 = (w10521 & ~w11361) | (w10521 & w18243) | (~w11361 & w18243);
assign w17337 = (w10531 & ~w10826) | (w10531 & w18244) | (~w10826 & w18244);
assign w17338 = (w10548 & ~w11117) | (w10548 & w18245) | (~w11117 & w18245);
assign w17339 = (w10517 & ~w11020) | (w10517 & w18246) | (~w11020 & w18246);
assign w17340 = (w10546 & ~w10964) | (w10546 & w18247) | (~w10964 & w18247);
assign w17341 = ~w11202 & w10523;
assign w17342 = (w10577 & ~w11020) | (w10577 & w18248) | (~w11020 & w18248);
assign w17343 = (w10585 & ~w11361) | (w10585 & w18249) | (~w11361 & w18249);
assign w17344 = ~w11245 & w10583;
assign w17345 = (w10582 & ~w10964) | (w10582 & w18250) | (~w10964 & w18250);
assign w17346 = (w10581 & ~w11117) | (w10581 & w18251) | (~w11117 & w18251);
assign w17347 = (w10579 & ~w10826) | (w10579 & w18252) | (~w10826 & w18252);
assign w17348 = ~w11202 & w10571;
assign w17349 = ~w10052 & w10256;
assign w17350 = w1699 & w10545;
assign w17351 = w1699 & w16717;
assign w17352 = ~w3449 & w10576;
assign w17353 = ~w3449 & w16720;
assign w17354 = ~w2784 & w10578;
assign w17355 = ~w2784 & w16719;
assign w17356 = w11480 & w18253;
assign w17357 = w10064 & ~w10130;
assign w17358 = w10064 & w16726;
assign w17359 = ~w11202 & w10970;
assign w17360 = (w10967 & ~w11117) | (w10967 & w18254) | (~w11117 & w18254);
assign w17361 = ~w16624 & w4808;
assign w17362 = (w10861 & ~w11099) | (w10861 & w18255) | (~w11099 & w18255);
assign w17363 = ~w16624 & w4797;
assign w17364 = (w10891 & ~w11318) | (w10891 & w18256) | (~w11318 & w18256);
assign w17365 = w10549 & w2198;
assign w17366 = ~w11202 & w10865;
assign w17367 = (w10869 & ~w11117) | (w10869 & w18257) | (~w11117 & w18257);
assign w17368 = (w10868 & ~w10964) | (w10868 & w18258) | (~w10964 & w18258);
assign w17369 = ~w11245 & w10870;
assign w17370 = (w10871 & ~w11406) | (w10871 & w18259) | (~w11406 & w18259);
assign w17371 = w11912 & ~w9434;
assign w17372 = (~w10042 & w17371) | (~w10042 & w18260) | (w17371 & w18260);
assign w17373 = w11931 & w18261;
assign w17374 = ~w11319 & w11006;
assign w17375 = ~w10052 & w9955;
assign w17376 = (w11007 & ~w11406) | (w11007 & w18262) | (~w11406 & w18262);
assign w17377 = w9929 & ~w10130;
assign w17378 = w9929 & w16726;
assign w17379 = w7785 & ~w10130;
assign w17380 = w7785 & w16726;
assign w17381 = ~w10853 & w7787;
assign w17382 = w12001 & ~w7789;
assign w17383 = w12001 & ~w16752;
assign w17384 = w12002 & w18263;
assign w17385 = ~w984 & w10545;
assign w17386 = ~w984 & w16717;
assign w17387 = ~w311 & w10572;
assign w17388 = ~w311 & w16718;
assign w17389 = (w6266 & ~w10826) | (w6266 & w18264) | (~w10826 & w18264);
assign w17390 = ~w6265 & w12011;
assign w17391 = ~w11245 & w10817;
assign w17392 = ~w11042 & w10836;
assign w17393 = w12067 & w18265;
assign w17394 = (w11176 & ~w11384) | (w11176 & w18266) | (~w11384 & w18266);
assign w17395 = ~w11245 & w11162;
assign w17396 = ~w1043 & w10545;
assign w17397 = ~w1043 & w16717;
assign w17398 = (w11169 & ~w11318) | (w11169 & w18267) | (~w11318 & w18267);
assign w17399 = ~w11168 & w12108;
assign w17400 = w12088 & w18268;
assign w17401 = ~w12123 & ~pi012;
assign w17402 = ~w11407 & w11059;
assign w17403 = ~w11385 & w11069;
assign w17404 = ~w11245 & w11053;
assign w17405 = w12184 & ~pi011;
assign w17406 = ~w10601 & w11121;
assign w17407 = (w11109 & ~w10826) | (w11109 & w18269) | (~w10826 & w18269);
assign w17408 = ~w11202 & w11119;
assign w17409 = ~w11493 & w11111;
assign w17410 = ~w11365 & w11107;
assign w17411 = w12222 & ~w11123;
assign w17412 = w12222 & ~w16771;
assign w17413 = w10574 & ~w2291;
assign w17414 = ~w1104 & w10545;
assign w17415 = ~w1104 & w16717;
assign w17416 = (w11150 & ~w10826) | (w11150 & w18270) | (~w10826 & w18270);
assign w17417 = (w11148 & ~w11020) | (w11148 & w18271) | (~w11020 & w18271);
assign w17418 = w10192 & ~w10130;
assign w17419 = w10192 & w16726;
assign w17420 = w12267 & ~pi016;
assign w17421 = ~w11270 & w12290;
assign w17422 = ~w10601 & w11342;
assign w17423 = w10549 & ~w8895;
assign w17424 = ~w10601 & w11422;
assign w17425 = ~w9672 & w12384;
assign w17426 = (w11396 & ~w10944) | (w11396 & w18272) | (~w10944 & w18272);
assign w17427 = w12418 & w12330;
assign w17428 = ~w1757 & ~w1230;
assign w17429 = ~w1757 & ~w1420;
assign w17430 = ~w1757 & w3331;
assign w17431 = ~w3346 & ~w1949;
assign w17432 = w342 & ~w2383;
assign w17433 = w342 & w16223;
assign w17434 = w16831 & w5424;
assign w17435 = (w5424 & w16831) | (w5424 & w4853) | (w16831 & w4853);
assign w17436 = ~w4691 & w4788;
assign w17437 = w4848 & w5594;
assign w17438 = ~w2723 & ~w5504;
assign w17439 = w6354 & ~w3949;
assign w17440 = ~w6390 & w6098;
assign w17441 = ~w6390 & w5224;
assign w17442 = w6305 & ~w5481;
assign w17443 = ~w6390 & w3683;
assign w17444 = ~w6390 & ~w4519;
assign w17445 = ~w6390 & w2695;
assign w17446 = w6224 & w6204;
assign w17447 = ~w6390 & w2444;
assign w17448 = ~w6390 & ~w7119;
assign w17449 = ~w6141 & ~w7148;
assign w17450 = ~w6552 & w7165;
assign w17451 = ~w6411 & w7194;
assign w17452 = ~w6552 & w7115;
assign w17453 = ~w6411 & w7119;
assign w17454 = ~w6411 & w7148;
assign w17455 = ~w6552 & ~w6219;
assign w17456 = ~w6552 & w6422;
assign w17457 = w6427 & w6473;
assign w17458 = ~w6411 & w6476;
assign w17459 = ~w6552 & w6469;
assign w17460 = ~w6552 & w6524;
assign w17461 = ~w6411 & w6545;
assign w17462 = ~w6411 & w6611;
assign w17463 = ~w6411 & w6560;
assign w17464 = w6427 & w6581;
assign w17465 = ~w6552 & w6568;
assign w17466 = w7882 & w7966;
assign w17467 = ~w8049 & w8031;
assign w17468 = ~w7806 & w9632;
assign w17469 = w16878 | w9183;
assign w17470 = (w9183 & w16878) | (w9183 & ~w9395) | (w16878 & ~w9395);
assign w17471 = ~w7806 & w9030;
assign w17472 = ~w7806 & w9213;
assign w17473 = ~w7806 & w9184;
assign w17474 = ~w7806 & w9991;
assign w17475 = ~w7806 & w9448;
assign w17476 = ~w7806 & w9489;
assign w17477 = ~w7806 & w9115;
assign w17478 = ~w7806 & w9149;
assign w17479 = w10212 & w9701;
assign w17480 = w5494 & ~w5529;
assign w17481 = w4841 & w3405;
assign w17482 = ~w1292 & w4009;
assign w17483 = ~w1292 & w5452;
assign w17484 = ~w1292 & ~w4163;
assign w17485 = ~w1292 & ~w4313;
assign w17486 = ~w1292 & ~w2753;
assign w17487 = ~w17029 & w4696;
assign w17488 = ~w3980 & w4695;
assign w17489 = ~w3980 & w4793;
assign w17490 = ~w17029 & w4789;
assign w17491 = ~w3980 & w4833;
assign w17492 = w6175 & w6162;
assign w17493 = ~w3743 & w5424;
assign w17494 = w6175 & w6221;
assign w17495 = w6175 & w6237;
assign w17496 = w6175 & w6303;
assign w17497 = w6175 & w6143;
assign w17498 = ~w6556 & w3019;
assign w17499 = ~w6529 & w6500;
assign w17500 = ~w6556 & ~w2990;
assign w17501 = ~w6556 & w6241;
assign w17502 = ~w6529 & w6640;
assign w17503 = w7684 & w7176;
assign w17504 = ~w7206 & w7168;
assign w17505 = w7684 & w7225;
assign w17506 = w7684 & w7175;
assign w17507 = w7684 & w7632;
assign w17508 = ~w7206 & ~w7113;
assign w17509 = w7684 & w7651;
assign w17510 = ~w7206 & w7655;
assign w17511 = ~w7206 & w7813;
assign w17512 = w7684 & w7808;
assign w17513 = w7684 & w7756;
assign w17514 = w7684 & w7868;
assign w17515 = ~w7206 & w7829;
assign w17516 = w7684 & w7841;
assign w17517 = (w9044 & ~w8463) | (w9044 & w17938) | (~w8463 & w17938);
assign w17518 = (w8417 & ~w8463) | (w8417 & w17939) | (~w8463 & w17939);
assign w17519 = (w8360 & ~w8463) | (w8360 & w17940) | (~w8463 & w17940);
assign w17520 = w8348 & w7980;
assign w17521 = (w7970 & ~w8463) | (w7970 & w17941) | (~w8463 & w17941);
assign w17522 = (w8345 & ~w8463) | (w8345 & w17942) | (~w8463 & w17942);
assign w17523 = w8347 & w18273;
assign w17524 = (w8441 & ~w8463) | (w8441 & w17943) | (~w8463 & w17943);
assign w17525 = w8348 & w8472;
assign w17526 = (w8597 & ~w8463) | (w8597 & w17944) | (~w8463 & w17944);
assign w17527 = w8348 & w8594;
assign w17528 = (w8526 & ~w8463) | (w8526 & w17945) | (~w8463 & w17945);
assign w17529 = w8348 & w8517;
assign w17530 = w8348 & w8573;
assign w17531 = (w8634 & ~w8463) | (w8634 & w17946) | (~w8463 & w17946);
assign w17532 = w8348 & w8680;
assign w17533 = ~w3295 & w3400;
assign w17534 = ~w3437 & w3440;
assign w17535 = ~w3465 & w3468;
assign w17536 = ~w3496 & w3497;
assign w17537 = ~w3522 & w3525;
assign w17538 = w3603 & ~pi180;
assign w17539 = ~w3603 & pi180;
assign w17540 = w3752 & ~pi260;
assign w17541 = ~w3752 & pi260;
assign w17542 = w3783 & ~w3782;
assign w17543 = w3839 & ~pi252;
assign w17544 = ~w3839 & pi252;
assign w17545 = w3870 & ~w3869;
assign w17546 = w2539 & ~w2502;
assign w17547 = ~w3405 & w3351;
assign w17548 = w3391 & ~w1292;
assign w17549 = ~w3405 & w4075;
assign w17550 = ~w3401 & w4076;
assign w17551 = ~w3401 & w3357;
assign w17552 = ~w4830 & w4769;
assign w17553 = ~w4830 & w4770;
assign w17554 = ~w4756 & w4771;
assign w17555 = (w4777 & w4832) | (w4777 & w17947) | (w4832 & w17947);
assign w17556 = ~w4099 & ~w3352;
assign w17557 = w16254 & w3920;
assign w17558 = (w3920 & w16254) | (w3920 & w4099) | (w16254 & w4099);
assign w17559 = ~w4756 & w5436;
assign w17560 = ~w5426 & w16255;
assign w17561 = w3391 & ~w1104;
assign w17562 = ~w3405 & w3350;
assign w17563 = ~w4853 & w5476;
assign w17564 = w16257 & w5478;
assign w17565 = (w5478 & w16257) | (w5478 & w4853) | (w16257 & w4853);
assign w17566 = w4677 & w2229;
assign w17567 = w16260 & w5513;
assign w17568 = (w5513 & w16260) | (w5513 & w4099) | (w16260 & w4099);
assign w17569 = w17053 & w5529;
assign w17570 = ~w4830 & w4832;
assign w17571 = ~w5593 & w4839;
assign w17572 = w16268 | ~w4687;
assign w17573 = (~w4687 & w16268) | (~w4687 & ~w5459) | (w16268 & ~w5459);
assign w17574 = ~w5638 & ~w5637;
assign w17575 = w4774 & ~w2695;
assign w17576 = ~w6208 & w6201;
assign w17577 = ~w6208 & w16291;
assign w17578 = (w5415 & ~w5597) | (w5415 & w18101) | (~w5597 & w18101);
assign w17579 = (w5415 & w16294) | (w5415 & ~w5608) | (w16294 & ~w5608);
assign w17580 = w6227 & w6230;
assign w17581 = ~w5530 & w5522;
assign w17582 = ~w5555 & ~w4831;
assign w17583 = w6286 & w6293;
assign w17584 = ~w6222 & ~w6296;
assign w17585 = w16320 & w6322;
assign w17586 = (w6322 & w16320) | (w6322 & w5480) | (w16320 & w5480);
assign w17587 = w6144 & w6379;
assign w17588 = ~w6169 & w6396;
assign w17589 = ~w16324 & w6404;
assign w17590 = ~w6169 & w6425;
assign w17591 = ~w16324 & w6154;
assign w17592 = w6305 & w6431;
assign w17593 = ~w6169 & w5629;
assign w17594 = ~w16324 & w5637;
assign w17595 = ~w16324 & w6471;
assign w17596 = ~w16324 & w6288;
assign w17597 = ~w6169 & w6275;
assign w17598 = (w6291 & ~w6177) | (w6291 & w17948) | (~w6177 & w17948);
assign w17599 = ~w16324 & w6224;
assign w17600 = ~w6169 & w6208;
assign w17601 = ~w16324 & w6197;
assign w17602 = ~w6545 & w17949;
assign w17603 = w6549 & ~w16351;
assign w17604 = ~w16324 & w6175;
assign w17605 = w6145 & w2564;
assign w17606 = ~w5643 & w6173;
assign w17607 = w5598 & ~w5461;
assign w17608 = ~w6293 & w17607;
assign w17609 = ~w6169 & ~w5407;
assign w17610 = ~w16324 & w6236;
assign w17611 = ~w6169 & w6249;
assign w17612 = ~w2164 & w6614;
assign w17613 = ~w16324 & w6321;
assign w17614 = ~w6305 & w6314;
assign w17615 = ~w6169 & w6312;
assign w17616 = ~w6261 & w6300;
assign w17617 = ~w16324 & w6302;
assign w17618 = w7105 & w7112;
assign w17619 = ~w16324 & w6174;
assign w17620 = ~w16324 & w7137;
assign w17621 = ~w6329 & w6380;
assign w17622 = (w6963 & ~w7151) | (w6963 & w18102) | (~w7151 & w18102);
assign w17623 = ~w883 & w7146;
assign w17624 = (~w883 & ~w6585) | (~w883 & w18103) | (~w6585 & w18103);
assign w17625 = ~w6553 & w6455;
assign w17626 = w17158 & w17950;
assign w17627 = ~w5341 & w6580;
assign w17628 = ~w5341 & w16372;
assign w17629 = ~w7191 & w7614;
assign w17630 = w249 & w7146;
assign w17631 = (w249 & ~w6585) | (w249 & w18274) | (~w6585 & w18274);
assign w17632 = w4371 & ~w16345;
assign w17633 = ~w6446 & w7633;
assign w17634 = (w6397 & ~w6438) | (w6397 & w18275) | (~w6438 & w18275);
assign w17635 = ~w6553 & w6410;
assign w17636 = ~w6446 & ~w5828;
assign w17637 = ~w7655 & ~w6412;
assign w17638 = ~w7655 & w6461;
assign w17639 = ~w7191 & w5857;
assign w17640 = (w7699 & w6494) | (w7699 & w17951) | (w6494 & w17951);
assign w17641 = ~w7191 & ~w4400;
assign w17642 = ~w7171 & w6677;
assign w17643 = ~w2229 & ~w5431;
assign w17644 = (w3623 & ~w7151) | (w3623 & w18104) | (~w7151 & w18104);
assign w17645 = w723 & w7146;
assign w17646 = w723 & ~w7182;
assign w17647 = w3197 & w6580;
assign w17648 = w3197 & w16372;
assign w17649 = ~w6627 & w6543;
assign w17650 = ~w3048 & w6412;
assign w17651 = ~w3048 & ~w6461;
assign w17652 = (w2723 & ~w7151) | (w2723 & w18105) | (~w7151 & w18105);
assign w17653 = ~w6553 & w7815;
assign w17654 = w2291 & w6412;
assign w17655 = w2291 & ~w6461;
assign w17656 = (w659 & ~w7151) | (w659 & w18106) | (~w7151 & w18106);
assign w17657 = ~w6553 & w6650;
assign w17658 = ~w6627 & w6641;
assign w17659 = (w1137 & ~w7151) | (w1137 & w18276) | (~w7151 & w18276);
assign w17660 = ~w6446 & w6631;
assign w17661 = ~w7906 & w18277;
assign w17662 = w7911 & w6461;
assign w17663 = w1670 & ~w6639;
assign w17664 = w1670 & ~w16411;
assign w17665 = (w7195 & ~w7669) | (w7195 & w17952) | (~w7669 & w17952);
assign w17666 = w7926 & w7958;
assign w17667 = (w7174 & ~w17666) | (w7174 & w17953) | (~w17666 & w17953);
assign w17668 = ~w7628 & w6999;
assign w17669 = (w7188 & ~w7837) | (w7188 & w18107) | (~w7837 & w18107);
assign w17670 = ~w7898 & w7223;
assign w17671 = ~w7959 & w7224;
assign w17672 = (w7222 & ~w7837) | (w7222 & w18108) | (~w7837 & w18108);
assign w17673 = (~w6447 & ~w7669) | (~w6447 & w18278) | (~w7669 & w18278);
assign w17674 = (w7639 & ~w7837) | (w7639 & w18279) | (~w7837 & w18279);
assign w17675 = (w7629 & ~w7711) | (w7629 & w17954) | (~w7711 & w17954);
assign w17676 = ~w7628 & ~w8369;
assign w17677 = (w7609 & ~w17666) | (w7609 & w17955) | (~w17666 & w17955);
assign w17678 = (w7610 & ~w7711) | (w7610 & w17956) | (~w7711 & w17956);
assign w17679 = ~w7628 & ~w7565;
assign w17680 = (w8408 & ~w7669) | (w8408 & w17957) | (~w7669 & w17957);
assign w17681 = (w8412 & ~w17666) | (w8412 & w17958) | (~w17666 & w17958);
assign w17682 = ~w3225 & w7166;
assign w17683 = (~w3225 & ~w7804) | (~w3225 & w17959) | (~w7804 & w17959);
assign w17684 = ~w7700 & w8437;
assign w17685 = (w7665 & ~w7837) | (w7665 & w18109) | (~w7837 & w18109);
assign w17686 = ~w7628 & ~w5769;
assign w17687 = ~w7782 & w7667;
assign w17688 = (w7664 & ~w17666) | (w7664 & w17960) | (~w17666 & w17960);
assign w17689 = w8437 & w18491;
assign w17690 = (w7705 & ~w7791) | (w7705 & w18280) | (~w7791 & w18280);
assign w17691 = (w7743 & ~w17666) | (w7743 & w18281) | (~w17666 & w18281);
assign w17692 = (w7801 & ~w7669) | (w7801 & w17961) | (~w7669 & w17961);
assign w17693 = (~w8556 & ~w7628) | (~w8556 & w17962) | (~w7628 & w17962);
assign w17694 = (w7809 & ~w7837) | (w7809 & w18111) | (~w7837 & w18111);
assign w17695 = ~w7814 & ~w8558;
assign w17696 = (w7799 & ~w17666) | (w7799 & w17963) | (~w17666 & w17963);
assign w17697 = (w7760 & ~w7669) | (w7760 & w17964) | (~w7669 & w17964);
assign w17698 = ~w7628 & ~w3565;
assign w17699 = (w7755 & ~w17666) | (w7755 & w17965) | (~w17666 & w17965);
assign w17700 = w6307 & ~w7759;
assign w17701 = (w7763 & ~w7837) | (w7763 & w18112) | (~w7837 & w18112);
assign w17702 = ~w7628 & ~w249;
assign w17703 = (w7867 & ~w7837) | (w7867 & w18113) | (~w7837 & w18113);
assign w17704 = (w7864 & ~w17666) | (w7864 & w17966) | (~w17666 & w17966);
assign w17705 = (w7861 & ~w7669) | (w7861 & w17967) | (~w7669 & w17967);
assign w17706 = (w7840 & ~w17666) | (w7840 & w17968) | (~w17666 & w17968);
assign w17707 = ~w8697 & w7844;
assign w17708 = (w7839 & ~w7837) | (w7839 & w18114) | (~w7837 & w18114);
assign w17709 = ~w7628 & ~w2322;
assign w17710 = ~w8378 & ~w7648;
assign w17711 = ~w8378 & w8406;
assign w17712 = (w7982 & ~w8429) | (w7982 & w18115) | (~w8429 & w18115);
assign w17713 = ~w8378 & w7964;
assign w17714 = ~w8378 & w8443;
assign w17715 = (w8435 & ~w8429) | (w8435 & w18116) | (~w8429 & w18116);
assign w17716 = w9261 & w9264;
assign w17717 = (w8610 & ~w17255) | (w8610 & w18282) | (~w17255 & w18282);
assign w17718 = w9305 & w8593;
assign w17719 = ~w8378 & w8527;
assign w17720 = ~w8430 & w8558;
assign w17721 = ~w8378 & w8630;
assign w17722 = ~w8430 & w8660;
assign w17723 = ~w8430 & w7993;
assign w17724 = ~w9110 & w9009;
assign w17725 = (w9642 & ~w17718) | (w9642 & w17969) | (~w17718 & w17969);
assign w17726 = ~w9265 & w9644;
assign w17727 = (w9346 & ~w9339) | (w9346 & w17970) | (~w9339 & w17970);
assign w17728 = (w9554 & ~w9339) | (w9554 & w17971) | (~w9339 & w17971);
assign w17729 = ~w9056 & w9545;
assign w17730 = (w9555 & ~w9447) | (w9555 & w17972) | (~w9447 & w17972);
assign w17731 = (w9553 & ~w17716) | (w9553 & w17973) | (~w17716 & w17973);
assign w17732 = (w9045 & ~w17716) | (w9045 & w17974) | (~w17716 & w17974);
assign w17733 = (w9028 & ~w17718) | (w9028 & w17975) | (~w17718 & w17975);
assign w17734 = (w9041 & ~w9339) | (w9041 & w17976) | (~w9339 & w17976);
assign w17735 = (w9048 & ~w9447) | (w9048 & w17977) | (~w9447 & w17977);
assign w17736 = ~w9307 & w9064;
assign w17737 = ~w9362 & w9073;
assign w17738 = ~w9473 & w9072;
assign w17739 = ~w9476 & w9065;
assign w17740 = ~w9056 & w9070;
assign w17741 = (w9068 & ~w17716) | (w9068 & w17978) | (~w17716 & w17978);
assign w17742 = ~w9110 & w9067;
assign w17743 = ~w9110 & w9210;
assign w17744 = (w9212 & ~w17718) | (w9212 & w17979) | (~w17718 & w17979);
assign w17745 = (w9224 & ~w17716) | (w9224 & w17980) | (~w17716 & w17980);
assign w17746 = ~w9056 & w9201;
assign w17747 = ~w9179 & w9116;
assign w17748 = (w9186 & ~w9447) | (w9186 & w17981) | (~w9447 & w17981);
assign w17749 = (w9187 & ~w9339) | (w9187 & w17982) | (~w9339 & w17982);
assign w17750 = (w9189 & ~w17716) | (w9189 & w17983) | (~w17716 & w17983);
assign w17751 = (w9188 & ~w17718) | (w9188 & w17984) | (~w17718 & w17984);
assign w17752 = ~w9056 & w9256;
assign w17753 = ~w9110 & w9248;
assign w17754 = (w9250 & ~w9178) | (w9250 & w17985) | (~w9178 & w17985);
assign w17755 = (~w8516 & ~w17716) | (~w8516 & w17986) | (~w17716 & w17986);
assign w17756 = (w9348 & ~w9509) | (w9348 & w18462) | (~w9509 & w18462);
assign w17757 = (w9333 & ~w17716) | (w9333 & w17987) | (~w17716 & w17987);
assign w17758 = (w9942 & ~w17718) | (w9942 & w17988) | (~w17718 & w17988);
assign w17759 = (w9297 & ~w9339) | (w9297 & w17989) | (~w9339 & w17989);
assign w17760 = (w9279 & ~w9447) | (w9279 & w17990) | (~w9447 & w17990);
assign w17761 = (w9296 & ~w17716) | (w9296 & w17991) | (~w17716 & w17991);
assign w17762 = ~w9056 & w9368;
assign w17763 = ~w9179 & w9374;
assign w17764 = (w9392 & ~w9447) | (w9392 & w17992) | (~w9447 & w17992);
assign w17765 = (w9372 & ~w17718) | (w9372 & w17993) | (~w17718 & w17993);
assign w17766 = (w9370 & ~w17716) | (w9370 & w17994) | (~w17716 & w17994);
assign w17767 = w10001 & w17995;
assign w17768 = (w9406 & ~w9447) | (w9406 & w17996) | (~w9447 & w17996);
assign w17769 = (w9440 & ~w17716) | (w9440 & w17997) | (~w17716 & w17997);
assign w17770 = (w9450 & ~w17718) | (w9450 & w17998) | (~w17718 & w17998);
assign w17771 = ~w9056 & w9454;
assign w17772 = (w9507 & ~w9339) | (w9507 & w17999) | (~w9339 & w17999);
assign w17773 = (w9487 & ~w17718) | (w9487 & w18000) | (~w17718 & w18000);
assign w17774 = ~w9056 & w9478;
assign w17775 = ~w9473 & w9506;
assign w17776 = ~w9265 & w9483;
assign w17777 = ~w9179 & w9491;
assign w17778 = ~w9362 & w9125;
assign w17779 = ~w9056 & w9124;
assign w17780 = ~w9110 & w9120;
assign w17781 = ~w9265 & w9126;
assign w17782 = (w9127 & ~w9447) | (w9127 & w18001) | (~w9447 & w18001);
assign w17783 = (w9119 & ~w17718) | (w9119 & w18002) | (~w17718 & w18002);
assign w17784 = ~w9362 & w9145;
assign w17785 = ~w9473 & w9144;
assign w17786 = ~w7378 & w9660;
assign w17787 = ~w9781 & w17786;
assign w17788 = ~w10184 & w16581;
assign w17789 = ~w10119 & w10528;
assign w17790 = (w9656 & ~w9692) | (w9656 & w18003) | (~w9692 & w18003);
assign w17791 = ~w10119 & w10258;
assign w17792 = ~w10184 & w10248;
assign w17793 = (w10033 & ~w9692) | (w10033 & w18004) | (~w9692 & w18004);
assign w17794 = (w10121 & ~w10183) | (w10121 & w18283) | (~w10183 & w18283);
assign w17795 = (w10056 & ~w10183) | (w10056 & w18284) | (~w10183 & w18284);
assign w17796 = (w9937 & ~w10183) | (w9937 & w18285) | (~w10183 & w18285);
assign w17797 = ~w10119 & w9834;
assign w17798 = (w9859 & ~w9692) | (w9859 & w18005) | (~w9692 & w18005);
assign w17799 = ~w10184 & w9768;
assign w17800 = w10553 & ~w9701;
assign w17801 = w10553 & ~w16627;
assign w17802 = ~w10119 & w9759;
assign w17803 = (w10217 & ~w10183) | (w10217 & w18286) | (~w10183 & w18286);
assign w17804 = w9125 & ~w9363;
assign w17805 = (w9125 & ~w9921) | (w9125 & w18006) | (~w9921 & w18006);
assign w17806 = (w10177 & ~w9692) | (w10177 & w18007) | (~w9692 & w18007);
assign w17807 = (w11291 & ~w10183) | (w11291 & w18287) | (~w10183 & w18287);
assign w17808 = (w9704 & ~w9692) | (w9704 & w18008) | (~w9692 & w18008);
assign w17809 = ~w10119 & w9707;
assign w17810 = w16690 | w9703;
assign w17811 = (w9703 & w16690) | (w9703 & ~w10005) | (w16690 & ~w10005);
assign w17812 = (w9712 & ~w10183) | (w9712 & w18288) | (~w10183 & w18288);
assign w17813 = (w9733 & ~w10183) | (w9733 & w18289) | (~w10183 & w18289);
assign w17814 = ~w10184 & w9678;
assign w17815 = ~w10184 & w9655;
assign w17816 = (w10972 & ~w10620) | (w10972 & w18009) | (~w10620 & w18009);
assign w17817 = ~w1668 & w10512;
assign w17818 = (~w1668 & ~w11243) | (~w1668 & w18010) | (~w11243 & w18010);
assign w17819 = w10072 & ~w9730;
assign w17820 = (w10072 & ~w11362) | (w10072 & w18011) | (~w11362 & w18011);
assign w17821 = w11823 & w18012;
assign w17822 = (w10036 & ~w11362) | (w10036 & w18013) | (~w11362 & w18013);
assign w17823 = (w10860 & ~w10565) | (w10860 & w18014) | (~w10565 & w18014);
assign w17824 = (w11003 & ~w10565) | (w11003 & w18015) | (~w10565 & w18015);
assign w17825 = (~w12015 & ~w11990) | (~w12015 & w18016) | (~w11990 & w18016);
assign w17826 = (w11170 & ~w10565) | (w11170 & w18017) | (~w10565 & w18017);
assign w17827 = (w11164 & ~w10620) | (w11164 & w18018) | (~w10620 & w18018);
assign w17828 = w12206 & w18019;
assign w17829 = ~w12235 & ~w12251;
assign w17830 = w12306 & w12304;
assign w17831 = w12324 & w11476;
assign w17832 = ~w10627 & w11338;
assign w17833 = ~w10567 & w11343;
assign w17834 = w12349 & ~w9730;
assign w17835 = w12349 & ~w11364;
assign w17836 = w12363 & w12330;
assign w17837 = w7317 & w10512;
assign w17838 = (w7317 & ~w11243) | (w7317 & w18020) | (~w11243 & w18020);
assign w17839 = (w9628 & ~w11362) | (w9628 & w18021) | (~w11362 & w18021);
assign w17840 = w12208 & w18290;
assign w17841 = w5412 & w5600;
assign w17842 = w5412 & w5511;
assign w17843 = w5412 & w5413;
assign w17844 = w5412 & w5551;
assign w17845 = ~w9895 & w9708;
assign w17846 = ~w9895 & w9657;
assign w17847 = ~w11360 & w11024;
assign w17848 = w4775 & ~w4071;
assign w17849 = w4775 & w4745;
assign w17850 = w4775 & w4698;
assign w17851 = w4775 & w4794;
assign w17852 = ~w5479 & ~w5629;
assign w17853 = ~w5477 & ~w6135;
assign w17854 = ~w5479 & w883;
assign w17855 = w5506 | w16834;
assign w17856 = ~w5479 & ~w3048;
assign w17857 = w5552 | w16838;
assign w17858 = ~w5479 & w2291;
assign w17859 = w5633 & ~w5481;
assign w17860 = w5633 & w6279;
assign w17861 = w5633 & w6243;
assign w17862 = w5633 & w6311;
assign w17863 = w6676 & ~w6307;
assign w17864 = w6452 & w6412;
assign w17865 = ~w6575 & w7147;
assign w17866 = ~w6575 & w6673;
assign w17867 = ~w7880 & w7185;
assign w17868 = ~w7880 & w7613;
assign w17869 = ~w7880 & w8410;
assign w17870 = ~w7600 & w6098;
assign w17871 = ~w7880 & w7652;
assign w17872 = ~w7880 & w7805;
assign w17873 = ~w7600 & w2695;
assign w17874 = w7600 & w8599;
assign w17875 = ~w7880 & w7776;
assign w17876 = ~w7819 & w7869;
assign w17877 = ~w7880 & w7847;
assign w17878 = ~w7600 & w2444;
assign w17879 = ~w7130 & ~w6392;
assign w17880 = ~w7130 & w6503;
assign w17881 = ~w7130 & w6488;
assign w17882 = ~w7130 & w16402;
assign w17883 = ~w7130 & w6579;
assign w17884 = (w7764 & ~w7217) | (w7764 & w18117) | (~w7217 & w18117);
assign w17885 = ~w7207 & w7766;
assign w17886 = ~w7218 & w7904;
assign w17887 = (w7907 & ~w7837) | (w7907 & w18291) | (~w7837 & w18291);
assign w17888 = ~w7823 & w7905;
assign w17889 = ~w7628 & w1168;
assign w17890 = ~w7884 & w7903;
assign w17891 = (w7922 & ~w7693) | (w7922 & w18292) | (~w7693 & w18292);
assign w17892 = ~w7959 & w8640;
assign w17893 = w8645 & ~w8632;
assign w17894 = ~w3949 & w821;
assign w17895 = ~w6180 & ~w4847;
assign w17896 = ~w7207 & w7860;
assign w17897 = ~w7218 & w7863;
assign w17898 = ~w7823 & w7843;
assign w17899 = ~w7700 & w7833;
assign w17900 = ~w7626 & ~w7993;
assign w17901 = w9014 & w7146;
assign w17902 = w9014 & ~w7182;
assign w17903 = ~w7761 & w5432;
assign w17904 = ~w8335 & w7979;
assign w17905 = ~w8318 & ~w7259;
assign w17906 = ~w8318 & w7057;
assign w17907 = ~w8515 & w16463;
assign w17908 = ~w8515 & w8327;
assign w17909 = (w8453 & ~w8399) | (w8453 & w18293) | (~w8399 & w18293);
assign w17910 = ~w8335 & w8528;
assign w17911 = (w8570 & ~w8323) | (w8570 & w18294) | (~w8323 & w18294);
assign w17912 = ~w6521 & w8561;
assign w17913 = ~w8335 & w8698;
assign w17914 = ~w8335 & w8625;
assign w17915 = w628 & w10572;
assign w17916 = w628 & w16718;
assign w17917 = ~w7988 & w8419;
assign w17918 = ~w7988 & w8392;
assign w17919 = ~w7988 & w8454;
assign w17920 = ~w7988 & w8482;
assign w17921 = w5475 & ~w4839;
assign w17922 = ~w17029 & w4676;
assign w17923 = ~w5477 & w16272;
assign w17924 = ~w5407 & w18492;
assign w17925 = w5438 & w6389;
assign w17926 = w6175 & w6346;
assign w17927 = w5633 & w6205;
assign w17928 = w6175 & w6198;
assign w17929 = ~w6575 & w7146;
assign w17930 = ~w17137 & w6452;
assign w17931 = ~w17137 & w7138;
assign w17932 = w6452 & w6423;
assign w17933 = ~w17137 & w6678;
assign w17934 = ~w6529 & w6544;
assign w17935 = w6676 & w6601;
assign w17936 = ~w6529 & w6567;
assign w17937 = ~w6575 & w6632;
assign w17938 = w5431 & w9044;
assign w17939 = w5431 & w8417;
assign w17940 = w5431 & w8360;
assign w17941 = w5431 & w7970;
assign w17942 = w5431 & w8345;
assign w17943 = w5431 & w8441;
assign w17944 = w5431 & w8597;
assign w17945 = w5431 & w8526;
assign w17946 = w5431 & w8634;
assign w17947 = ~w17029 & w4777;
assign w17948 = w6175 & w6291;
assign w17949 = w6202 & ~w6204;
assign w17950 = w7150 & w7583;
assign w17951 = ~w6405 & w7699;
assign w17952 = ~w17640 & w7195;
assign w17953 = ~w7927 & w7174;
assign w17954 = ~w7752 & w7629;
assign w17955 = ~w7927 & w7609;
assign w17956 = ~w7752 & w7610;
assign w17957 = ~w17640 & w8408;
assign w17958 = ~w7927 & w8412;
assign w17959 = (~w3225 & w7805) | (~w3225 & w18295) | (w7805 & w18295);
assign w17960 = ~w7927 & w7664;
assign w17961 = ~w17640 & w7801;
assign w17962 = ~w2932 & ~w8556;
assign w17963 = ~w7927 & w7799;
assign w17964 = ~w17640 & w7760;
assign w17965 = ~w7927 & w7755;
assign w17966 = ~w7927 & w7864;
assign w17967 = ~w17640 & w7861;
assign w17968 = ~w7927 & w7840;
assign w17969 = ~w9304 & w9642;
assign w17970 = ~w9361 & w9346;
assign w17971 = (w9554 & ~w9331) | (w9554 & w18296) | (~w9331 & w18296);
assign w17972 = (w9555 & ~w9439) | (w9555 & w18297) | (~w9439 & w18297);
assign w17973 = ~w9262 & w9553;
assign w17974 = (w9045 & ~w9259) | (w9045 & w18298) | (~w9259 & w18298);
assign w17975 = ~w9304 & w9028;
assign w17976 = ~w9361 & w9041;
assign w17977 = ~w9472 & w9048;
assign w17978 = ~w9262 & w9068;
assign w17979 = ~w9304 & w9212;
assign w17980 = ~w9262 & w9224;
assign w17981 = (w9186 & ~w9439) | (w9186 & w18299) | (~w9439 & w18299);
assign w17982 = (w9187 & ~w9331) | (w9187 & w18300) | (~w9331 & w18300);
assign w17983 = (w9189 & ~w9259) | (w9189 & w18463) | (~w9259 & w18463);
assign w17984 = (w9188 & ~w9303) | (w9188 & w18301) | (~w9303 & w18301);
assign w17985 = w9172 & w9250;
assign w17986 = ~w9262 & ~w8516;
assign w17987 = (w9333 & ~w9259) | (w9333 & w18302) | (~w9259 & w18302);
assign w17988 = ~w9304 & w9942;
assign w17989 = ~w9361 & w9297;
assign w17990 = ~w9472 & w9279;
assign w17991 = ~w9262 & w9296;
assign w17992 = (w9392 & ~w9439) | (w9392 & w18303) | (~w9439 & w18303);
assign w17993 = (w9372 & ~w9303) | (w9372 & w18304) | (~w9303 & w18304);
assign w17994 = ~w9262 & w9370;
assign w17995 = w10002 & w10007;
assign w17996 = (w9406 & ~w9439) | (w9406 & w18305) | (~w9439 & w18305);
assign w17997 = ~w9262 & w9440;
assign w17998 = ~w9304 & w9450;
assign w17999 = ~w9361 & w9507;
assign w18000 = ~w9304 & w9487;
assign w18001 = ~w9472 & w9127;
assign w18002 = ~w9304 & w9119;
assign w18003 = ~w9693 & w9656;
assign w18004 = ~w9693 & w10033;
assign w18005 = ~w9693 & w9859;
assign w18006 = (w9125 & w9901) | (w9125 & w18306) | (w9901 & w18306);
assign w18007 = ~w9693 & w10177;
assign w18008 = ~w9693 & w9704;
assign w18009 = ~w16607 & w10972;
assign w18010 = ~w11242 & ~w1668;
assign w18011 = ~w11363 & w10072;
assign w18012 = ~w11812 & w18307;
assign w18013 = ~w11363 & w10036;
assign w18014 = ~w10566 & w10860;
assign w18015 = ~w10566 & w11003;
assign w18016 = ~w11989 & ~w12015;
assign w18017 = ~w10566 & w11170;
assign w18018 = ~w16607 & w11164;
assign w18019 = ~w12200 & ~w5889;
assign w18020 = ~w11242 & w7317;
assign w18021 = ~w11363 & w9628;
assign w18022 = ~w4756 & ~w4051;
assign w18023 = ~w5530 & w5537;
assign w18024 = ~w5538 & w5533;
assign w18025 = w6276 & w18308;
assign w18026 = w6281 & ~w16295;
assign w18027 = w6284 & w6286;
assign w18028 = ~w6169 & w6340;
assign w18029 = ~w6305 & w6342;
assign w18030 = w6145 & w1388;
assign w18031 = ~w17073 & w2873;
assign w18032 = ~w6305 & w6203;
assign w18033 = ~w6169 & w6181;
assign w18034 = ~w17073 & ~w6098;
assign w18035 = ~w17073 & ~w5857;
assign w18036 = ~w1073 & ~w6649;
assign w18037 = ~w6178 & w6561;
assign w18038 = ~w7134 & w7189;
assign w18039 = ~w2291 & ~w6607;
assign w18040 = ~w6516 & w7116;
assign w18041 = ~w1358 & ~w6649;
assign w18042 = w2416 & ~w6607;
assign w18043 = ~w17618 & ~w6963;
assign w18044 = w7134 & ~w6557;
assign w18045 = ~w1168 & w6382;
assign w18046 = ~w1168 & ~w6649;
assign w18047 = w2322 & w6406;
assign w18048 = w2322 & ~w6607;
assign w18049 = w7645 & w7628;
assign w18050 = ~w7130 & w6393;
assign w18051 = ~w7130 & w6424;
assign w18052 = ~w6493 & w6497;
assign w18053 = w2753 & w7165;
assign w18054 = w2753 & ~w6557;
assign w18055 = ~w6446 & w6506;
assign w18056 = ~w7766 & ~w6473;
assign w18057 = ~w7766 & ~w16394;
assign w18058 = ~w17618 & w2961;
assign w18059 = ~w6596 & ~w4797;
assign w18060 = ~w7130 & w6599;
assign w18061 = ~w7130 & w6633;
assign w18062 = (w7214 & ~w7217) | (w7214 & w18309) | (~w7217 & w18309);
assign w18063 = (w7630 & ~w7205) | (w7630 & w18310) | (~w7205 & w18310);
assign w18064 = ~w7207 & w7606;
assign w18065 = ~w7823 & w7608;
assign w18066 = w5192 & w7175;
assign w18067 = w5192 & w17207;
assign w18068 = ~w7087 & ~w7113;
assign w18069 = ~w7087 & w17213;
assign w18070 = (w7674 & ~w7217) | (w7674 & w18311) | (~w7217 & w18311);
assign w18071 = (w7703 & ~w7205) | (w7703 & w18312) | (~w7205 & w18312);
assign w18072 = ~w7823 & w7717;
assign w18073 = (w7714 & ~w7837) | (w7714 & w18313) | (~w7837 & w18313);
assign w18074 = (w7720 & ~w7693) | (w7720 & w18314) | (~w7693 & w18314);
assign w18075 = ~w7218 & w7810;
assign w18076 = w7806 & w8556;
assign w18077 = w7806 & ~w17693;
assign w18078 = (w9978 & ~w9664) | (w9978 & w18464) | (~w9664 & w18464);
assign w18079 = (w10036 & ~w9727) | (w10036 & w18315) | (~w9727 & w18315);
assign w18080 = (w10105 & ~w9664) | (w10105 & w18465) | (~w9664 & w18465);
assign w18081 = (w10100 & ~w9727) | (w10100 & w18316) | (~w9727 & w18316);
assign w18082 = (w9952 & ~w9727) | (w9952 & w18317) | (~w9727 & w18317);
assign w18083 = (w9938 & ~w9664) | (w9938 & w18466) | (~w9664 & w18466);
assign w18084 = (w9815 & ~w9664) | (w9815 & w18467) | (~w9664 & w18467);
assign w18085 = (w9844 & ~w9727) | (w9844 & w18318) | (~w9727 & w18318);
assign w18086 = (w10153 & ~w9727) | (w10153 & w18319) | (~w9727 & w18319);
assign w18087 = (w9702 & ~w9664) | (w9702 & w18468) | (~w9664 & w18468);
assign w18088 = ~w9728 & w9628;
assign w18089 = ~w9665 & w11427;
assign w18090 = w7591 & w7164;
assign w18091 = w7591 & w7683;
assign w18092 = w7591 & w7762;
assign w18093 = w7591 & w7866;
assign w18094 = ~w9961 & w9643;
assign w18095 = w5449 | w16840;
assign w18096 = w6175 & w6398;
assign w18097 = w6175 & w5646;
assign w18098 = w6175 & w16368;
assign w18099 = ~w8397 & w8368;
assign w18100 = ~w8397 & w7983;
assign w18101 = w5415 | w16835;
assign w18102 = ~w7190 & w6963;
assign w18103 = ~w7181 & ~w883;
assign w18104 = ~w7190 & w3623;
assign w18105 = ~w7190 & w2723;
assign w18106 = ~w7190 & w659;
assign w18107 = ~w17193 & w7188;
assign w18108 = ~w17193 & w7222;
assign w18109 = ~w17193 & w7665;
assign w18110 = w7698 & ~w7663;
assign w18111 = ~w17193 & w7809;
assign w18112 = ~w17193 & w7763;
assign w18113 = ~w17193 & w7867;
assign w18114 = ~w17193 & w7839;
assign w18115 = ~w8428 & w7982;
assign w18116 = ~w8428 & w8435;
assign w18117 = w7215 & w7764;
assign w18118 = w16302 | w5550;
assign w18119 = (w5550 & w16302) | (w5550 & ~w5538) | (w16302 & ~w5538);
assign w18120 = w11984 & w11991;
assign w18121 = ~w12004 & pi009;
assign w18122 = w9973 & ~w11364;
assign w18123 = w11000 & ~w3048;
assign w18124 = ~w10567 & w10832;
assign w18125 = ~w10627 & w10838;
assign w18126 = ~w11319 & w10813;
assign w18127 = ~w11100 & w10830;
assign w18128 = w4924 & w10520;
assign w18129 = w4924 & ~w11364;
assign w18130 = ~w10601 & w11171;
assign w18131 = ~w11319 & w11054;
assign w18132 = w9891 & ~w11364;
assign w18133 = ~w10627 & w11079;
assign w18134 = ~w12186 & ~w12137;
assign w18135 = ~w10567 & w11285;
assign w18136 = ~w11464 & ~w11478;
assign w18137 = w7259 & w10512;
assign w18138 = w7259 & ~w11244;
assign w18139 = ~w10627 & w17423;
assign w18140 = ~w10567 & w11423;
assign w18141 = w7347 & w10512;
assign w18142 = w7347 & ~w11244;
assign w18143 = ~w10567 & w11218;
assign w18144 = w10549 & ~w7288;
assign w18145 = w9766 & ~w9730;
assign w18146 = w9766 & ~w11364;
assign w18147 = w12444 & w10512;
assign w18148 = w12444 & ~w11244;
assign w18149 = w12458 & ~pi019;
assign w18150 = ~w12458 & ~pi018;
assign w18151 = w12418 & w16818;
assign w18152 = w12363 & w16821;
assign w18153 = w12424 & ~w16131;
assign w18154 = w12424 & ~w16148;
assign w18155 = w5860 & w5481;
assign w18156 = w7591 & w7910;
assign w18157 = ~w8499 & ~w4580;
assign w18158 = w9555 & w9032;
assign w18159 = w9555 & w9123;
assign w18160 = ~w9895 & w10525;
assign w18161 = ~w9895 & ~w9363;
assign w18162 = ~w9895 & w10253;
assign w18163 = w10212 & w9979;
assign w18164 = w10841 & ~w9975;
assign w18165 = ~w9895 & w10019;
assign w18166 = w9741 & w10010;
assign w18167 = ~w8462 & w10032;
assign w18168 = w10212 & w10011;
assign w18169 = w10127 & w16895;
assign w18170 = ~w8462 & w10060;
assign w18171 = ~w16559 & w9955;
assign w18172 = ~w9438 & w9953;
assign w18173 = w9171 & w11047;
assign w18174 = w10212 & w9910;
assign w18175 = ~w16559 & w9885;
assign w18176 = w10212 & w9795;
assign w18177 = ~w9895 & w9830;
assign w18178 = ~w9895 & w9856;
assign w18179 = ~w9438 & w9878;
assign w18180 = w10212 & w9849;
assign w18181 = w9741 & w9847;
assign w18182 = ~w9895 & w9758;
assign w18183 = ~w16559 & w10211;
assign w18184 = ~w9895 & w10213;
assign w18185 = ~w8462 & w10212;
assign w18186 = ~w16559 & w10160;
assign w18187 = w10212 & w10155;
assign w18188 = w9741 & w10154;
assign w18189 = ~w8462 & w10158;
assign w18190 = ~w9438 & w10178;
assign w18191 = ~w9971 & w9703;
assign w18192 = ~w9895 & w9732;
assign w18193 = ~w16559 & w9735;
assign w18194 = ~w8462 & w9736;
assign w18195 = ~w9438 & w9739;
assign w18196 = ~w11360 & w10520;
assign w18197 = ~w11360 & ~w9730;
assign w18198 = ~w11360 & w10910;
assign w18199 = w11374 & w10932;
assign w18200 = ~w16649 & w10913;
assign w18201 = ~w16612 & w10911;
assign w18202 = ~w9899 & w11031;
assign w18203 = ~w10988 & w11023;
assign w18204 = ~w16649 & w11009;
assign w18205 = ~w16612 & w11029;
assign w18206 = ~w11360 & w11278;
assign w18207 = ~w11360 & w11390;
assign w18208 = ~w16612 & w11389;
assign w18209 = ~w9899 & w11223;
assign w18210 = ~w10988 & w11221;
assign w18211 = w11374 & w11212;
assign w18212 = ~w16649 & w11226;
assign w18213 = ~w9931 & w11219;
assign w18214 = ~w16612 & w11220;
assign w18215 = ~w9422 & w10050;
assign w18216 = w9634 & w17266;
assign w18217 = w9634 & w16533;
assign w18218 = ~w16881 & ~w9434;
assign w18219 = ~w9799 & ~w5889;
assign w18220 = ~w16881 & w9711;
assign w18221 = ~w16899 & w10580;
assign w18222 = ~w16893 & w10578;
assign w18223 = ~w16893 & w10951;
assign w18224 = ~w16893 & w10866;
assign w18225 = w5769 & w10857;
assign w18226 = ~w16893 & w11196;
assign w18227 = ~w16899 & w11271;
assign w18228 = ~w16893 & w11275;
assign w18229 = ~w16893 & w11340;
assign w18230 = ~w16899 & w11412;
assign w18231 = ~w16893 & w11418;
assign w18232 = ~w5479 & w4163;
assign w18233 = ~w17137 & w6569;
assign w18234 = ~w17137 & w6637;
assign w18235 = w6452 & w6643;
assign w18236 = ~w8397 & w8681;
assign w18237 = ~w8499 & ~w9634;
assign w18238 = ~w17301 & w10897;
assign w18239 = w10176 & ~w17312;
assign w18240 = w10176 & ~w17313;
assign w18241 = ~w9438 & w10190;
assign w18242 = w11098 & w10552;
assign w18243 = ~w11360 & w10521;
assign w18244 = ~w16612 & w10531;
assign w18245 = ~w16649 & w10548;
assign w18246 = ~w9931 & w10517;
assign w18247 = ~w10988 & w10546;
assign w18248 = ~w9931 & w10577;
assign w18249 = ~w11360 & w10585;
assign w18250 = ~w10988 & w10582;
assign w18251 = ~w16649 & w10581;
assign w18252 = ~w16612 & w10579;
assign w18253 = w11761 & pi024;
assign w18254 = ~w16649 & w10967;
assign w18255 = w11098 & w10861;
assign w18256 = w11312 & w10891;
assign w18257 = ~w16649 & w10869;
assign w18258 = ~w10988 & w10868;
assign w18259 = w11399 & w10871;
assign w18260 = w11912 & w16894;
assign w18261 = w11932 & pi005;
assign w18262 = w11399 & w11007;
assign w18263 = ~w11997 & ~pi010;
assign w18264 = ~w16612 & w6266;
assign w18265 = w12068 & pi007;
assign w18266 = w11374 & w11176;
assign w18267 = w11312 & w11169;
assign w18268 = ~w12081 & w8462;
assign w18269 = ~w16612 & w11109;
assign w18270 = ~w16612 & w11150;
assign w18271 = ~w9931 & w11148;
assign w18272 = ~w9015 & w11396;
assign w18273 = w691 & w8440;
assign w18274 = ~w7181 & w249;
assign w18275 = w6427 & w6397;
assign w18276 = ~w7190 & w1137;
assign w18277 = ~w1168 & ~w6643;
assign w18278 = ~w17640 & ~w6447;
assign w18279 = ~w17193 & w7639;
assign w18280 = ~w7790 & w7705;
assign w18281 = ~w7927 & w7743;
assign w18282 = ~w8387 & w8610;
assign w18283 = ~w10176 & w10121;
assign w18284 = ~w10176 & w10056;
assign w18285 = ~w10176 & w9937;
assign w18286 = ~w10176 & w10217;
assign w18287 = ~w10176 & w11291;
assign w18288 = ~w10176 & w9712;
assign w18289 = ~w10176 & w9733;
assign w18290 = w17828 & pi015;
assign w18291 = ~w17193 & w7907;
assign w18292 = w7684 & w7922;
assign w18293 = ~w8397 & w8453;
assign w18294 = w8325 & w8570;
assign w18295 = ~w7824 & ~w3225;
assign w18296 = ~w16489 & w9554;
assign w18297 = ~w1699 & w9555;
assign w18298 = w9251 & w9045;
assign w18299 = ~w1699 & w9186;
assign w18300 = ~w16489 & w9187;
assign w18301 = ~w9302 & w9188;
assign w18302 = w9251 & w9333;
assign w18303 = ~w1699 & w9392;
assign w18304 = ~w9302 & w9372;
assign w18305 = ~w1699 & w9406;
assign w18306 = ~w9899 & w9125;
assign w18307 = ~w11811 & pi003;
assign w18308 = ~w6275 & ~w5413;
assign w18309 = w7215 & w7214;
assign w18310 = ~w7206 & w7630;
assign w18311 = w7215 & w7674;
assign w18312 = ~w7206 & w7703;
assign w18313 = ~w17193 & w7714;
assign w18314 = w7684 & w7720;
assign w18315 = ~w9718 & w10036;
assign w18316 = ~w9718 & w10100;
assign w18317 = ~w9718 & w9952;
assign w18318 = ~w9718 & w9844;
assign w18319 = ~w9718 & w10153;
assign w18320 = w4684 & ~w4104;
assign w18321 = ~w5480 & w1104;
assign w18322 = ~w6178 & w6319;
assign w18323 = ~w6178 & w5645;
assign w18324 = ~w6493 & w7118;
assign w18325 = ~w6516 & w6428;
assign w18326 = ~w7706 & w7752;
assign w18327 = w1388 & ~w6649;
assign w18328 = ~w17618 & w1073;
assign w18329 = w6377 & ~w6649;
assign w18330 = w7645 & ~w7626;
assign w18331 = ~w7753 & w7588;
assign w18332 = ~w7782 & w7677;
assign w18333 = w7173 & ~w1043;
assign w18334 = ~w7898 & w7682;
assign w18335 = ~w7207 & w7678;
assign w18336 = ~w7898 & w7740;
assign w18337 = w6307 & w7704;
assign w18338 = ~w7823 & w7761;
assign w18339 = ~w7207 & w7906;
assign w18340 = w8637 & ~w6649;
assign w18341 = ~w8430 & w9077;
assign w18342 = ~w8430 & w8529;
assign w18343 = ~w8378 & w8716;
assign w18344 = ~w7967 & w9481;
assign w18345 = ~w8378 & w8659;
assign w18346 = w16519 | ~w8051;
assign w18347 = (~w8051 & w16519) | (~w8051 & ~w9562) | (w16519 & ~w9562);
assign w18348 = ~w9473 & w9222;
assign w18349 = ~w9088 & w16520;
assign w18350 = ~w9088 & w9549;
assign w18351 = ~w9362 & w9101;
assign w18352 = ~w9088 & w9094;
assign w18353 = ~w9265 & w9099;
assign w18354 = ~w9473 & w16532;
assign w18355 = ~w9088 & ~w8432;
assign w18356 = w9782 & w9781;
assign w18357 = ~w9088 & w9225;
assign w18358 = w9873 & w9881;
assign w18359 = w16546 | w9342;
assign w18360 = (w9342 & w16546) | (w9342 & ~w9562) | (w16546 & ~w9562);
assign w18361 = ~w9088 & w9330;
assign w18362 = ~w9056 & w9341;
assign w18363 = ~w9307 & ~w9027;
assign w18364 = ~w9317 & w9327;
assign w18365 = ~w9110 & w9340;
assign w18366 = ~w9179 & w9343;
assign w18367 = ~w9088 & w9375;
assign w18368 = ~w9110 & w16553;
assign w18369 = ~w9362 & w9393;
assign w18370 = ~w7805 & w9971;
assign w18371 = ~w9110 & w9415;
assign w18372 = ~w9088 & w9403;
assign w18373 = ~w9179 & w16557;
assign w18374 = ~w9476 & w9400;
assign w18375 = ~w9307 & w9416;
assign w18376 = ~w9265 & w9407;
assign w18377 = ~w9433 & w10038;
assign w18378 = w10089 & pi003;
assign w18379 = ~w9088 & w9117;
assign w18380 = ~w9362 & w9164;
assign w18381 = ~w9307 & w9170;
assign w18382 = ~w9473 & w9168;
assign w18383 = ~w10251 & w10250;
assign w18384 = ~w9307 & w17283;
assign w18385 = ~w9647 & w17284;
assign w18386 = ~w9265 & w17285;
assign w18387 = ~w9473 & w17286;
assign w18388 = w10267 & w10272;
assign w18389 = w16591 | w9634;
assign w18390 = (w9634 & w16591) | (w9634 & ~w9747) | (w16591 & ~w9747);
assign w18391 = ~w9926 & w9831;
assign w18392 = ~w10119 & w9682;
assign w18393 = ~w10184 & w16597;
assign w18394 = w17296 & w10810;
assign w18395 = (w10810 & w17296) | (w10810 & w10119) | (w17296 & w10119);
assign w18396 = ~w10184 & w9972;
assign w18397 = ~w10184 & w16615;
assign w18398 = ~w9825 & w10097;
assign w18399 = ~w9696 & w10092;
assign w18400 = ~w10226 & w10073;
assign w18401 = ~w10119 & w10064;
assign w18402 = ~w9696 & w10066;
assign w18403 = ~w9696 & w9954;
assign w18404 = ~w10226 & w9932;
assign w18405 = w11016 & w9931;
assign w18406 = ~w10119 & w9887;
assign w18407 = ~w9825 & w9906;
assign w18408 = ~w10089 & w9890;
assign w18409 = ~w10184 & w9907;
assign w18410 = w11064 & w9899;
assign w18411 = ~w10184 & w9793;
assign w18412 = ~w9696 & w9798;
assign w18413 = ~w9825 & w11132;
assign w18414 = ~w10184 & w16657;
assign w18415 = ~w10119 & w9848;
assign w18416 = ~w9696 & w16662;
assign w18417 = ~w11227 & ~w11228;
assign w18418 = ~w10119 & w10218;
assign w18419 = ~w10089 & w10214;
assign w18420 = ~w10119 & w10192;
assign w18421 = ~w11319 & w10812;
assign w18422 = ~w11158 & w11000;
assign w18423 = ~w10567 & ~w10532;
assign w18424 = ~w4687 & w11507;
assign w18425 = ~w7407 & w10512;
assign w18426 = ~w7407 & ~w11244;
assign w18427 = ~w9672 & w10544;
assign w18428 = ~w7378 & w10512;
assign w18429 = ~w7378 & ~w11244;
assign w18430 = ~w11090 & w10526;
assign w18431 = ~w11090 & w10588;
assign w18432 = ~w10590 & w11724;
assign w18433 = w11728 & ~w11715;
assign w18434 = ~w11158 & w10954;
assign w18435 = ~w11158 & w10926;
assign w18436 = ~w11319 & w10925;
assign w18437 = ~w10567 & w10933;
assign w18438 = ~w9672 & w10105;
assign w18439 = ~w10627 & w17365;
assign w18440 = ~w11909 & ~w11910;
assign w18441 = w17399 & w12108;
assign w18442 = (w12108 & w17399) | (w12108 & w11158) | (w17399 & w11158);
assign w18443 = w12292 & w11475;
assign w18444 = ~w11090 & w11368;
assign w18445 = w12351 & ~w12333;
assign w18446 = ~w12463 & ~w12483;
assign w18447 = w12247 & pi014;
assign w18448 = ~w9646 & w9185;
assign w18449 = ~w9646 & w9417;
assign w18450 = ~w11240 & w10512;
assign w18451 = ~w11240 & w10906;
assign w18452 = w16931 | w10856;
assign w18453 = (w10856 & w16931) | (w10856 & ~w11064) | (w16931 & ~w11064);
assign w18454 = ~w11240 & w11028;
assign w18455 = ~w11240 & w11125;
assign w18456 = w16959 | w11151;
assign w18457 = (w11151 & w16959) | (w11151 & ~w11064) | (w16959 & ~w11064);
assign w18458 = w16964 | w11287;
assign w18459 = (w11287 & w16964) | (w11287 & ~w10962) | (w16964 & ~w10962);
assign w18460 = w16967 | w11276;
assign w18461 = (w11276 & w16967) | (w11276 & ~w11064) | (w16967 & ~w11064);
assign w18462 = ~w9646 & w9348;
assign w18463 = w9251 & w9189;
assign w18464 = w9659 & w9978;
assign w18465 = w9659 & w10105;
assign w18466 = w9659 & w9938;
assign w18467 = w9659 & w9815;
assign w18468 = w9659 & w9702;
assign w18469 = (~w7171 & ~w1073) | (~w7171 & w18036) | (~w1073 & w18036);
assign w18470 = (~w6627 & ~w2291) | (~w6627 & w18039) | (~w2291 & w18039);
assign w18471 = (~w7171 & ~w1358) | (~w7171 & w18041) | (~w1358 & w18041);
assign w18472 = (~w6627 & w2416) | (~w6627 & w18042) | (w2416 & w18042);
assign w18473 = (~w6516 & w4371) | (~w6516 & w17632) | (w4371 & w17632);
assign w18474 = (w4400 & w7145) | (w4400 & ~w17641) | (w7145 & ~w17641);
assign w18475 = (~w7171 & w1388) | (~w7171 & w18327) | (w1388 & w18327);
assign w18476 = (~w7171 & w6377) | (~w7171 & w18329) | (w6377 & w18329);
assign w18477 = (~w7171 & w8637) | (~w7171 & w18340) | (w8637 & w18340);
assign w18478 = w7626 | ~w7647;
assign w18479 = (~w7989 & ~w7028) | (~w7989 & w17264) | (~w7028 & w17264);
assign w18480 = (~w9647 & w7626) | (~w9647 & w17267) | (w7626 & w17267);
assign w18481 = (~w8051 & w16519) | (~w8051 & ~w9566) | (w16519 & ~w9566);
assign w18482 = (~w9647 & w7903) | (~w9647 & w17277) | (w7903 & w17277);
assign w18483 = (w10570 & w16715) | (w10570 & ~w11195) | (w16715 & ~w11195);
assign w18484 = (~w11256 & w11041) | (~w11256 & ~w16817) | (w11041 & ~w16817);
assign w18485 = (w5475 & w17921) | (w5475 & ~w5597) | (w17921 & ~w5597);
assign w18486 = w5345 & ~w5377;
assign w18487 = (w5494 & w17480) | (w5494 & ~w5523) | (w17480 & ~w5523);
assign w18488 = w18486 & w5345;
assign w18489 = w18155 & w5860;
assign w18490 = w6327 & w6318;
assign w18491 = (~w7700 & w7698) | (~w7700 & w18110) | (w7698 & w18110);
assign w18492 = (w5345 & w18486) | (w5345 & w5479) | (w18486 & w5479);
assign one = 1;
assign po000 = pi000;
assign po001 = ~w921;
assign po002 = ~w1766;
assign po003 = ~w2580;
assign po004 = ~w3344;
assign po005 = ~w4091;
assign po006 = ~w4866;
assign po007 = ~w5627;
assign po008 = ~w6374;
assign po009 = ~w7163;
assign po010 = ~w7956;
assign po011 = ~w8747;
assign po012 = ~w9626;
assign po013 = ~w10511;
assign po014 = w11462;
assign po015 = w12511;
assign po016 = pi031;
assign po017 = pi032;
assign po018 = pi033;
assign po019 = pi034;
assign po020 = pi035;
assign po021 = pi036;
assign po022 = pi037;
assign po023 = pi038;
assign po024 = w12519;
assign po025 = ~w12522;
assign po026 = ~w12525;
assign po027 = ~w12528;
assign po028 = ~w12531;
assign po029 = ~w12534;
assign po030 = ~w12537;
assign po031 = ~w12540;
assign po032 = ~w12549;
assign po033 = ~w12557;
assign po034 = ~w12565;
assign po035 = ~w12573;
assign po036 = ~w12581;
assign po037 = ~w12589;
assign po038 = ~w12597;
assign po039 = ~w12605;
assign po040 = ~w12620;
assign po041 = ~w12629;
assign po042 = ~w12638;
assign po043 = ~w12647;
assign po044 = ~w12656;
assign po045 = ~w12665;
assign po046 = ~w12674;
assign po047 = ~w12683;
assign po048 = ~w12704;
assign po049 = ~w12718;
assign po050 = ~w12732;
assign po051 = ~w12746;
assign po052 = ~w12760;
assign po053 = ~w12774;
assign po054 = ~w12788;
assign po055 = ~w12802;
assign po056 = ~w12828;
assign po057 = ~w12844;
assign po058 = ~w12860;
assign po059 = ~w12875;
assign po060 = ~w12891;
assign po061 = ~w12907;
assign po062 = ~w12923;
assign po063 = ~w12938;
assign po064 = ~w12964;
assign po065 = ~w12985;
assign po066 = ~w13005;
assign po067 = ~w13025;
assign po068 = ~w13045;
assign po069 = ~w13065;
assign po070 = ~w13085;
assign po071 = ~w13105;
assign po072 = ~w13149;
assign po073 = ~w13171;
assign po074 = ~w13193;
assign po075 = ~w13214;
assign po076 = ~w13236;
assign po077 = ~w13258;
assign po078 = ~w13279;
assign po079 = ~w13300;
assign po080 = ~w13336;
assign po081 = ~w13366;
assign po082 = ~w13394;
assign po083 = ~w13425;
assign po084 = ~w13453;
assign po085 = ~w13481;
assign po086 = ~w13509;
assign po087 = ~w13538;
assign po088 = ~w13584;
assign po089 = ~w13615;
assign po090 = ~w13644;
assign po091 = ~w13677;
assign po092 = ~w13705;
assign po093 = ~w13735;
assign po094 = ~w13763;
assign po095 = ~w13792;
assign po096 = ~w13835;
assign po097 = ~w13874;
assign po098 = ~w13908;
assign po099 = ~w13941;
assign po100 = ~w13975;
assign po101 = ~w14008;
assign po102 = ~w14044;
assign po103 = ~w14079;
assign po104 = ~w14139;
assign po105 = ~w14175;
assign po106 = ~w14210;
assign po107 = ~w14245;
assign po108 = ~w14280;
assign po109 = ~w14315;
assign po110 = ~w14350;
assign po111 = ~w14385;
assign po112 = ~w14429;
assign po113 = ~w14466;
assign po114 = ~w14503;
assign po115 = ~w14540;
assign po116 = ~w14577;
assign po117 = ~w14614;
assign po118 = ~w14651;
assign po119 = ~w14688;
assign po120 = ~w14784;
assign po121 = ~w14825;
assign po122 = ~w14866;
assign po123 = ~w14907;
assign po124 = ~w14948;
assign po125 = ~w14989;
assign po126 = ~w15030;
assign po127 = ~w15071;
assign po128 = ~w15132;
assign po129 = ~w15185;
assign po130 = ~w15238;
assign po131 = ~w15291;
assign po132 = ~w15344;
assign po133 = ~w15397;
assign po134 = ~w15450;
assign po135 = ~w15503;
assign po136 = ~w15562;
assign po137 = ~w15617;
assign po138 = ~w15672;
assign po139 = ~w15727;
assign po140 = ~w15782;
assign po141 = ~w15837;
assign po142 = ~w15892;
assign po143 = ~w15947;
assign po144 = w29;
assign po145 = w955;
assign po146 = ~w15948;
assign po147 = ~w15950;
assign po148 = ~w15951;
assign po149 = w2632;
assign po150 = ~w15954;
assign po151 = ~w15955;
assign po152 = ~w15957;
assign po153 = ~w15959;
assign po154 = ~w15961;
assign po155 = ~w15965;
assign po156 = ~w15968;
assign po157 = ~w15970;
assign po158 = ~w15976;
assign po159 = ~w15979;
assign po160 = ~w15981;
assign po161 = w6392;
assign po162 = ~w15988;
assign po163 = ~w15991;
assign po164 = ~w15993;
assign po165 = ~w15995;
assign po166 = ~w16000;
assign po167 = ~w16002;
assign po168 = ~w16005;
assign po169 = ~w16009;
assign po170 = ~w16014;
assign po171 = ~w16018;
assign po172 = ~w16021;
assign po173 = ~w16027;
assign po174 = ~w16031;
assign po175 = ~w16035;
assign po176 = ~w16039;
assign po177 = ~w16047;
assign po178 = ~w16061;
assign po179 = ~w16064;
assign po180 = ~w16069;
assign po181 = ~w16075;
assign po182 = ~w16081;
assign po183 = w16087;
assign po184 = ~w16097;
assign po185 = ~w16103;
assign po186 = ~w16110;
assign po187 = ~w16118;
assign po188 = ~w16129;
assign po189 = ~w16138;
assign po190 = ~w16145;
assign po191 = ~w16151;
assign po192 = ~w16167;
endmodule

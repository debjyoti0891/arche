module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095;
assign w0 = pi00 & pi32;
assign w1 = pi01 & pi32;
assign w2 = pi00 & pi33;
assign w3 = w1 & ~w2;
assign w4 = ~w1 & w2;
assign w5 = ~w3 & ~w4;
assign w6 = ~pi33 & ~pi34;
assign w7 = pi33 & pi34;
assign w8 = ~w6 & ~w7;
assign w9 = pi00 & w8;
assign w10 = ~pi00 & pi33;
assign w11 = ~w1 & w10;
assign w12 = ~w9 & ~w11;
assign w13 = pi02 & pi32;
assign w14 = pi01 & ~pi32;
assign w15 = pi33 & ~w13;
assign w16 = ~w14 & w15;
assign w17 = ~pi33 & w13;
assign w18 = ~w16 & ~w17;
assign w19 = w12 & ~w18;
assign w20 = ~w12 & w18;
assign w21 = ~w19 & ~w20;
assign w22 = (w11 & w16) | (w11 & w8060) | (w16 & w8060);
assign w23 = ~pi35 & w7;
assign w24 = pi35 & w6;
assign w25 = ~w23 & ~w24;
assign w26 = pi00 & ~w25;
assign w27 = pi01 & w8;
assign w28 = (pi35 & w26) | (pi35 & w8061) | (w26 & w8061);
assign w29 = ~w26 & w8062;
assign w30 = ~w28 & ~w29;
assign w31 = pi03 & pi32;
assign w32 = pi02 & ~pi32;
assign w33 = pi33 & ~w31;
assign w34 = ~w32 & w33;
assign w35 = ~pi33 & w31;
assign w36 = ~w34 & ~w35;
assign w37 = w30 & ~w36;
assign w38 = ~w30 & w36;
assign w39 = ~w37 & ~w38;
assign w40 = (pi35 & ~w8) | (pi35 & w8063) | (~w8 & w8063);
assign w41 = (~w40 & w18) | (~w40 & w8064) | (w18 & w8064);
assign w42 = w39 & ~w41;
assign w43 = ~w39 & w41;
assign w44 = ~w42 & ~w43;
assign w45 = ~w22 & ~w44;
assign w46 = w22 & w44;
assign w47 = ~w45 & ~w46;
assign w48 = (~w42 & ~w44) | (~w42 & w8065) | (~w44 & w8065);
assign w49 = pi01 & ~w25;
assign w50 = pi02 & w8;
assign w51 = (pi35 & w49) | (pi35 & w7455) | (w49 & w7455);
assign w52 = ~w49 & w7456;
assign w53 = ~w51 & ~w52;
assign w54 = ~pi35 & ~pi36;
assign w55 = pi35 & pi36;
assign w56 = ~w54 & ~w55;
assign w57 = (pi37 & ~w56) | (pi37 & w7458) | (~w56 & w7458);
assign w58 = w56 & w8066;
assign w59 = ~w57 & ~w58;
assign w60 = w53 & ~w59;
assign w61 = ~w53 & w59;
assign w62 = ~w60 & ~w61;
assign w63 = pi04 & pi32;
assign w64 = pi03 & ~pi32;
assign w65 = pi33 & ~w63;
assign w66 = ~w64 & w65;
assign w67 = ~pi33 & w63;
assign w68 = ~w66 & ~w67;
assign w69 = w62 & ~w68;
assign w70 = ~w62 & w68;
assign w71 = ~w69 & ~w70;
assign w72 = w30 & w8067;
assign w73 = (~pi37 & ~w30) | (~pi37 & w8068) | (~w30 & w8068);
assign w74 = ~w72 & ~w73;
assign w75 = ~w71 & ~w74;
assign w76 = w71 & w74;
assign w77 = ~w75 & ~w76;
assign w78 = ~w48 & w77;
assign w79 = w48 & ~w77;
assign w80 = ~w78 & ~w79;
assign w81 = (~w60 & ~w62) | (~w60 & w8069) | (~w62 & w8069);
assign w82 = pi03 & w8;
assign w83 = (pi35 & ~w6) | (pi35 & w7457) | (~w6 & w7457);
assign w84 = w7 & w8070;
assign w85 = ~w82 & w8071;
assign w86 = pi35 & w82;
assign w87 = ~w85 & ~w86;
assign w88 = pi01 & w56;
assign w89 = (pi37 & ~w54) | (pi37 & w7458) | (~w54 & w7458);
assign w90 = ~pi37 & w55;
assign w91 = w55 & w8066;
assign w92 = ~w88 & w8072;
assign w93 = pi37 & w88;
assign w94 = ~w92 & ~w93;
assign w95 = w87 & w94;
assign w96 = ~w87 & ~w94;
assign w97 = ~w95 & ~w96;
assign w98 = pi05 & pi32;
assign w99 = pi04 & ~pi32;
assign w100 = pi33 & ~w98;
assign w101 = ~w99 & w100;
assign w102 = ~pi33 & w98;
assign w103 = ~w101 & ~w102;
assign w104 = w97 & ~w103;
assign w105 = ~w97 & w103;
assign w106 = ~w104 & ~w105;
assign w107 = ~w81 & w106;
assign w108 = w81 & ~w106;
assign w109 = ~w107 & ~w108;
assign w110 = (~w72 & ~w71) | (~w72 & w8073) | (~w71 & w8073);
assign w111 = w109 & ~w110;
assign w112 = ~w109 & w110;
assign w113 = ~w111 & ~w112;
assign w114 = ~w78 & ~w113;
assign w115 = w78 & w113;
assign w116 = ~w114 & ~w115;
assign w117 = ~pi37 & ~pi38;
assign w118 = pi37 & pi38;
assign w119 = ~w117 & ~w118;
assign w120 = pi00 & w119;
assign w121 = ~w95 & w103;
assign w122 = ~w121 & w7459;
assign w123 = (~w120 & w121) | (~w120 & w7460) | (w121 & w7460);
assign w124 = ~w122 & ~w123;
assign w125 = pi04 & w8;
assign w126 = (pi35 & ~w6) | (pi35 & w7461) | (~w6 & w7461);
assign w127 = w7 & w8074;
assign w128 = ~w125 & w8075;
assign w129 = pi35 & w125;
assign w130 = ~w128 & ~w129;
assign w131 = pi02 & w56;
assign w132 = (pi37 & ~w54) | (pi37 & w7462) | (~w54 & w7462);
assign w133 = w55 & w8076;
assign w134 = ~w131 & w8077;
assign w135 = pi37 & w131;
assign w136 = ~w134 & ~w135;
assign w137 = w130 & w136;
assign w138 = ~w130 & ~w136;
assign w139 = ~w137 & ~w138;
assign w140 = pi06 & pi32;
assign w141 = pi05 & ~pi32;
assign w142 = pi33 & ~w140;
assign w143 = ~w141 & w142;
assign w144 = ~pi33 & w140;
assign w145 = ~w143 & ~w144;
assign w146 = w139 & ~w145;
assign w147 = ~w139 & w145;
assign w148 = ~w146 & ~w147;
assign w149 = w124 & w148;
assign w150 = ~w124 & ~w148;
assign w151 = ~w149 & ~w150;
assign w152 = ~w111 & w8078;
assign w153 = (w151 & w111) | (w151 & w334) | (w111 & w334);
assign w154 = ~w152 & ~w153;
assign w155 = ~w115 & ~w154;
assign w156 = w115 & w154;
assign w157 = ~w155 & ~w156;
assign w158 = (pi39 & ~w119) | (pi39 & w8079) | (~w119 & w8079);
assign w159 = ~w122 & ~w158;
assign w160 = ~w149 & w159;
assign w161 = ~w121 & w8080;
assign w162 = w148 & w161;
assign w163 = ~w160 & ~w162;
assign w164 = ~w138 & ~w145;
assign w165 = pi39 & w117;
assign w166 = ~pi39 & w118;
assign w167 = ~w165 & ~w166;
assign w168 = pi00 & ~w167;
assign w169 = pi01 & w119;
assign w170 = (pi39 & w168) | (pi39 & w7463) | (w168 & w7463);
assign w171 = ~w168 & w7464;
assign w172 = ~w170 & ~w171;
assign w173 = ~w137 & ~w172;
assign w174 = ~w164 & w173;
assign w175 = ~w137 & w145;
assign w176 = ~w138 & w172;
assign w177 = ~w175 & w176;
assign w178 = ~w174 & ~w177;
assign w179 = pi05 & w8;
assign w180 = (pi35 & ~w6) | (pi35 & w7465) | (~w6 & w7465);
assign w181 = w7 & w8081;
assign w182 = ~w179 & w8082;
assign w183 = pi35 & w179;
assign w184 = ~w182 & ~w183;
assign w185 = pi03 & w56;
assign w186 = (pi37 & ~w54) | (pi37 & w7466) | (~w54 & w7466);
assign w187 = w55 & w8083;
assign w188 = ~w185 & w8084;
assign w189 = pi37 & w185;
assign w190 = ~w188 & ~w189;
assign w191 = w184 & w190;
assign w192 = ~w184 & ~w190;
assign w193 = ~w191 & ~w192;
assign w194 = pi07 & pi32;
assign w195 = pi06 & ~pi32;
assign w196 = pi33 & ~w194;
assign w197 = ~w195 & w196;
assign w198 = ~pi33 & w194;
assign w199 = ~w197 & ~w198;
assign w200 = w193 & ~w199;
assign w201 = ~w193 & w199;
assign w202 = ~w200 & ~w201;
assign w203 = w178 & ~w202;
assign w204 = ~w178 & w202;
assign w205 = ~w203 & ~w204;
assign w206 = ~w163 & w205;
assign w207 = w163 & ~w205;
assign w208 = ~w206 & ~w207;
assign w209 = ~w156 & w8085;
assign w210 = (w208 & w156) | (w208 & w213) | (w156 & w213);
assign w211 = ~w209 & ~w210;
assign w212 = w156 & w208;
assign w213 = w153 & w208;
assign w214 = ~w174 & ~w203;
assign w215 = ~pi39 & ~pi40;
assign w216 = pi39 & pi40;
assign w217 = ~w215 & ~w216;
assign w218 = pi00 & w217;
assign w219 = pi01 & ~w167;
assign w220 = pi02 & w119;
assign w221 = (pi39 & w219) | (pi39 & w7467) | (w219 & w7467);
assign w222 = ~w219 & w7468;
assign w223 = ~w221 & ~w222;
assign w224 = w218 & w223;
assign w225 = ~w218 & ~w223;
assign w226 = ~w224 & ~w225;
assign w227 = ~w191 & w199;
assign w228 = ~w192 & ~w227;
assign w229 = w226 & w228;
assign w230 = ~w226 & ~w228;
assign w231 = ~w229 & ~w230;
assign w232 = pi06 & w8;
assign w233 = (pi35 & ~w6) | (pi35 & w7469) | (~w6 & w7469);
assign w234 = w7 & w8086;
assign w235 = ~w232 & w8087;
assign w236 = pi35 & w232;
assign w237 = ~w235 & ~w236;
assign w238 = pi04 & w56;
assign w239 = (pi37 & ~w54) | (pi37 & w7470) | (~w54 & w7470);
assign w240 = w55 & w8088;
assign w241 = ~w238 & w8089;
assign w242 = pi37 & w238;
assign w243 = ~w241 & ~w242;
assign w244 = w237 & w243;
assign w245 = ~w237 & ~w243;
assign w246 = ~w244 & ~w245;
assign w247 = pi08 & pi32;
assign w248 = pi07 & ~pi32;
assign w249 = pi33 & ~w247;
assign w250 = ~w248 & w249;
assign w251 = ~pi33 & w247;
assign w252 = ~w250 & ~w251;
assign w253 = w246 & ~w252;
assign w254 = ~w246 & w252;
assign w255 = ~w253 & ~w254;
assign w256 = w231 & ~w255;
assign w257 = ~w231 & w255;
assign w258 = ~w256 & ~w257;
assign w259 = w214 & ~w258;
assign w260 = ~w214 & w258;
assign w261 = ~w259 & ~w260;
assign w262 = ~w162 & w205;
assign w263 = ~w160 & ~w262;
assign w264 = ~w261 & ~w263;
assign w265 = w261 & w263;
assign w266 = ~w264 & ~w265;
assign w267 = ~w213 & ~w266;
assign w268 = w213 & w266;
assign w269 = ~w267 & ~w268;
assign w270 = ~w212 & ~w269;
assign w271 = w212 & w269;
assign w272 = ~w270 & ~w271;
assign w273 = (pi41 & ~w217) | (pi41 & w8090) | (~w217 & w8090);
assign w274 = (~w273 & ~w223) | (~w273 & w8091) | (~w223 & w8091);
assign w275 = ~w230 & w255;
assign w276 = ~w275 & w7471;
assign w277 = (~w274 & w275) | (~w274 & w7472) | (w275 & w7472);
assign w278 = ~w276 & ~w277;
assign w279 = pi07 & w8;
assign w280 = w7 & w7473;
assign w281 = (pi35 & ~w6) | (pi35 & w8092) | (~w6 & w8092);
assign w282 = ~w279 & w8093;
assign w283 = pi35 & w279;
assign w284 = pi09 & pi32;
assign w285 = pi08 & ~pi32;
assign w286 = pi33 & ~w284;
assign w287 = ~w285 & w286;
assign w288 = ~pi33 & w284;
assign w289 = ~w287 & ~w288;
assign w290 = ~w282 & w7474;
assign w291 = (w289 & w282) | (w289 & w7475) | (w282 & w7475);
assign w292 = ~w290 & ~w291;
assign w293 = pi05 & w56;
assign w294 = (pi37 & ~w54) | (pi37 & w8094) | (~w54 & w8094);
assign w295 = pi04 & w90;
assign w296 = ~w293 & ~w294;
assign w297 = w56 & w8095;
assign w298 = (~w297 & ~w296) | (~w297 & w8096) | (~w296 & w8096);
assign w299 = w292 & ~w298;
assign w300 = ~w292 & w298;
assign w301 = ~w299 & ~w300;
assign w302 = ~pi41 & w216;
assign w303 = pi41 & w215;
assign w304 = ~w302 & ~w303;
assign w305 = pi00 & ~w304;
assign w306 = pi01 & w217;
assign w307 = (pi41 & w305) | (pi41 & w7476) | (w305 & w7476);
assign w308 = ~w305 & w7477;
assign w309 = ~w307 & ~w308;
assign w310 = pi02 & ~w167;
assign w311 = pi03 & w119;
assign w312 = (pi39 & w310) | (pi39 & w7478) | (w310 & w7478);
assign w313 = ~w310 & w7479;
assign w314 = ~w312 & ~w313;
assign w315 = w309 & w314;
assign w316 = ~w309 & ~w314;
assign w317 = ~w315 & ~w316;
assign w318 = ~w244 & w252;
assign w319 = ~w245 & ~w318;
assign w320 = w317 & w319;
assign w321 = ~w317 & ~w319;
assign w322 = ~w320 & ~w321;
assign w323 = w301 & ~w322;
assign w324 = ~w301 & w322;
assign w325 = ~w323 & ~w324;
assign w326 = w278 & ~w325;
assign w327 = ~w278 & w325;
assign w328 = ~w326 & ~w327;
assign w329 = ~w260 & w263;
assign w330 = ~w259 & ~w329;
assign w331 = ~w328 & ~w330;
assign w332 = w328 & w330;
assign w333 = ~w331 & ~w332;
assign w334 = w107 & w151;
assign w335 = w208 & w334;
assign w336 = w266 & w335;
assign w337 = w333 & w336;
assign w338 = ~w268 & ~w333;
assign w339 = ~w337 & ~w338;
assign w340 = w268 & w333;
assign w341 = ~w271 & ~w340;
assign w342 = w339 & ~w341;
assign w343 = ~w271 & ~w339;
assign w344 = ~w342 & ~w343;
assign w345 = pi43 & w315;
assign w346 = ~pi43 & ~w315;
assign w347 = ~w345 & ~w346;
assign w348 = w301 & ~w320;
assign w349 = (~w347 & w348) | (~w347 & w7480) | (w348 & w7480);
assign w350 = ~w348 & w7481;
assign w351 = ~w349 & ~w350;
assign w352 = (~w291 & ~w292) | (~w291 & w8097) | (~w292 & w8097);
assign w353 = ~pi41 & ~pi42;
assign w354 = pi41 & pi42;
assign w355 = ~w353 & ~w354;
assign w356 = (pi43 & ~w355) | (pi43 & w7486) | (~w355 & w7486);
assign w357 = w355 & w8098;
assign w358 = ~w356 & ~w357;
assign w359 = pi02 & w217;
assign w360 = (pi41 & ~w215) | (pi41 & w7482) | (~w215 & w7482);
assign w361 = w216 & w8099;
assign w362 = ~w359 & w8100;
assign w363 = pi41 & w359;
assign w364 = ~w362 & ~w363;
assign w365 = ~w358 & w364;
assign w366 = w358 & ~w364;
assign w367 = ~w365 & ~w366;
assign w368 = pi03 & ~w167;
assign w369 = pi04 & w119;
assign w370 = (pi39 & w368) | (pi39 & w8101) | (w368 & w8101);
assign w371 = ~w368 & w8102;
assign w372 = ~w370 & ~w371;
assign w373 = w367 & ~w372;
assign w374 = ~w367 & w372;
assign w375 = ~w373 & ~w374;
assign w376 = pi08 & w8;
assign w377 = pi33 & ~pi35;
assign w378 = ~w6 & ~w377;
assign w379 = ~pi34 & ~pi35;
assign w380 = pi07 & ~w379;
assign w381 = ~w378 & w380;
assign w382 = ~w376 & ~w381;
assign w383 = pi35 & ~w382;
assign w384 = ~pi35 & w382;
assign w385 = ~w383 & ~w384;
assign w386 = pi37 & ~w55;
assign w387 = pi06 & w56;
assign w388 = pi05 & ~w56;
assign w389 = ~w387 & ~w388;
assign w390 = w386 & ~w389;
assign w391 = (~pi37 & ~w55) | (~pi37 & w8103) | (~w55 & w8103);
assign w392 = ~w387 & w391;
assign w393 = ~w390 & ~w392;
assign w394 = w385 & w393;
assign w395 = ~w385 & ~w393;
assign w396 = ~w394 & ~w395;
assign w397 = pi10 & pi32;
assign w398 = pi09 & ~pi32;
assign w399 = pi33 & ~w397;
assign w400 = ~w398 & w399;
assign w401 = ~pi33 & w397;
assign w402 = ~w400 & ~w401;
assign w403 = w396 & ~w402;
assign w404 = ~w396 & w402;
assign w405 = ~w403 & ~w404;
assign w406 = w375 & ~w405;
assign w407 = ~w375 & w405;
assign w408 = ~w406 & ~w407;
assign w409 = w352 & w408;
assign w410 = ~w352 & ~w408;
assign w411 = ~w409 & ~w410;
assign w412 = ~w351 & ~w411;
assign w413 = w351 & w411;
assign w414 = ~w412 & ~w413;
assign w415 = ~w276 & ~w326;
assign w416 = ~w414 & ~w415;
assign w417 = w414 & w415;
assign w418 = ~w416 & ~w417;
assign w419 = (w418 & w337) | (w418 & w7483) | (w337 & w7483);
assign w420 = ~w337 & w7484;
assign w421 = ~w419 & ~w420;
assign w422 = ~w342 & ~w421;
assign w423 = w342 & w421;
assign w424 = ~w422 & ~w423;
assign w425 = pi04 & ~w167;
assign w426 = pi05 & w119;
assign w427 = (pi39 & w425) | (pi39 & w8104) | (w425 & w8104);
assign w428 = ~w425 & w8105;
assign w429 = ~w427 & ~w428;
assign w430 = pi03 & w217;
assign w431 = (pi41 & ~w215) | (pi41 & w7485) | (~w215 & w7485);
assign w432 = w216 & w8106;
assign w433 = ~w430 & w8107;
assign w434 = pi41 & w430;
assign w435 = ~w433 & ~w434;
assign w436 = pi01 & w355;
assign w437 = (pi43 & ~w353) | (pi43 & w7486) | (~w353 & w7486);
assign w438 = pi42 & ~pi43;
assign w439 = pi41 & w438;
assign w440 = w438 & w8108;
assign w441 = ~w436 & w8109;
assign w442 = pi43 & w436;
assign w443 = ~w441 & ~w442;
assign w444 = w435 & w443;
assign w445 = ~w435 & ~w443;
assign w446 = ~w444 & ~w445;
assign w447 = w429 & w446;
assign w448 = ~w429 & ~w446;
assign w449 = ~w447 & ~w448;
assign w450 = (~w394 & ~w396) | (~w394 & w7487) | (~w396 & w7487);
assign w451 = w449 & ~w450;
assign w452 = ~w449 & w450;
assign w453 = ~w451 & ~w452;
assign w454 = pi07 & w56;
assign w455 = (pi37 & ~w54) | (pi37 & w7488) | (~w54 & w7488);
assign w456 = w55 & w8110;
assign w457 = ~w454 & w8111;
assign w458 = pi37 & w454;
assign w459 = ~w457 & ~w458;
assign w460 = pi09 & w8;
assign w461 = (pi35 & ~w6) | (pi35 & w7489) | (~w6 & w7489);
assign w462 = w7 & w8112;
assign w463 = ~w460 & w8113;
assign w464 = pi35 & w460;
assign w465 = ~w463 & ~w464;
assign w466 = w459 & w465;
assign w467 = ~w459 & ~w465;
assign w468 = ~w466 & ~w467;
assign w469 = pi11 & pi32;
assign w470 = pi10 & ~pi32;
assign w471 = pi33 & ~w469;
assign w472 = ~w470 & w471;
assign w473 = ~pi33 & w469;
assign w474 = ~w472 & ~w473;
assign w475 = w468 & ~w474;
assign w476 = ~w468 & w474;
assign w477 = ~w475 & ~w476;
assign w478 = w453 & w477;
assign w479 = ~w453 & ~w477;
assign w480 = ~w478 & ~w479;
assign w481 = (~w366 & ~w367) | (~w366 & w8114) | (~w367 & w8114);
assign w482 = w408 & w7490;
assign w483 = (~w366 & ~w405) | (~w366 & w8115) | (~w405 & w8115);
assign w484 = (~w481 & w405) | (~w481 & w8116) | (w405 & w8116);
assign w485 = ~w483 & ~w484;
assign w486 = ~w352 & ~w481;
assign w487 = (w486 & ~w405) | (w486 & w8117) | (~w405 & w8117);
assign w488 = ~w485 & ~w487;
assign w489 = ~w482 & w488;
assign w490 = w480 & ~w489;
assign w491 = ~w480 & w489;
assign w492 = ~w490 & ~w491;
assign w493 = w411 & w7491;
assign w494 = ~w345 & ~w350;
assign w495 = (w494 & ~w411) | (w494 & w7492) | (~w411 & w7492);
assign w496 = ~w493 & ~w495;
assign w497 = w492 & ~w496;
assign w498 = ~w492 & w496;
assign w499 = ~w497 & ~w498;
assign w500 = w259 & ~w328;
assign w501 = (~w500 & ~w414) | (~w500 & w8118) | (~w414 & w8118);
assign w502 = ~w416 & ~w501;
assign w503 = w499 & w502;
assign w504 = ~w499 & ~w502;
assign w505 = ~w503 & ~w504;
assign w506 = w337 & w418;
assign w507 = w505 & w506;
assign w508 = w265 & ~w328;
assign w509 = w418 & w508;
assign w510 = w505 & w509;
assign w511 = ~w505 & ~w509;
assign w512 = ~w510 & ~w511;
assign w513 = w423 & w512;
assign w514 = ~w423 & ~w506;
assign w515 = ~w512 & w514;
assign w516 = ~w507 & ~w513;
assign w517 = ~w515 & w516;
assign w518 = (~w493 & w492) | (~w493 & w7871) | (w492 & w7871);
assign w519 = (~w481 & w485) | (~w481 & w8119) | (w485 & w8119);
assign w520 = (~w519 & ~w489) | (~w519 & w8120) | (~w489 & w8120);
assign w521 = ~pi43 & ~pi44;
assign w522 = pi43 & pi44;
assign w523 = ~w521 & ~w522;
assign w524 = pi00 & w523;
assign w525 = (~w444 & ~w446) | (~w444 & w8121) | (~w446 & w8121);
assign w526 = ~w524 & w525;
assign w527 = w524 & ~w525;
assign w528 = ~w526 & ~w527;
assign w529 = (~w451 & ~w453) | (~w451 & w7493) | (~w453 & w7493);
assign w530 = ~w528 & w529;
assign w531 = w528 & ~w529;
assign w532 = ~w530 & ~w531;
assign w533 = (~w466 & ~w468) | (~w466 & w7494) | (~w468 & w7494);
assign w534 = pi05 & ~w167;
assign w535 = pi06 & w119;
assign w536 = (pi39 & w534) | (pi39 & w8122) | (w534 & w8122);
assign w537 = ~w534 & w8123;
assign w538 = ~w536 & ~w537;
assign w539 = pi02 & w355;
assign w540 = (pi43 & ~w353) | (pi43 & w7495) | (~w353 & w7495);
assign w541 = w438 & w8124;
assign w542 = ~w539 & w8125;
assign w543 = pi43 & w539;
assign w544 = ~w542 & ~w543;
assign w545 = pi04 & w217;
assign w546 = (pi41 & ~w215) | (pi41 & w7496) | (~w215 & w7496);
assign w547 = w216 & w8126;
assign w548 = ~w545 & w8127;
assign w549 = pi41 & w545;
assign w550 = ~w548 & ~w549;
assign w551 = ~w544 & ~w550;
assign w552 = w544 & w550;
assign w553 = ~w551 & ~w552;
assign w554 = ~w538 & w553;
assign w555 = w538 & ~w553;
assign w556 = ~w554 & ~w555;
assign w557 = ~w533 & ~w556;
assign w558 = w533 & w556;
assign w559 = ~w557 & ~w558;
assign w560 = pi08 & w56;
assign w561 = (pi37 & ~w54) | (pi37 & w7497) | (~w54 & w7497);
assign w562 = w55 & w8128;
assign w563 = ~w560 & w8129;
assign w564 = pi37 & w560;
assign w565 = ~w563 & ~w564;
assign w566 = pi10 & w8;
assign w567 = (pi35 & ~w6) | (pi35 & w7498) | (~w6 & w7498);
assign w568 = w7 & w8130;
assign w569 = ~w566 & w8131;
assign w570 = pi35 & w566;
assign w571 = ~w569 & ~w570;
assign w572 = w565 & w571;
assign w573 = ~w565 & ~w571;
assign w574 = ~w572 & ~w573;
assign w575 = pi12 & pi32;
assign w576 = pi11 & ~pi32;
assign w577 = pi33 & ~w575;
assign w578 = ~w576 & w577;
assign w579 = ~pi33 & w575;
assign w580 = ~w578 & ~w579;
assign w581 = w574 & ~w580;
assign w582 = ~w574 & w580;
assign w583 = ~w581 & ~w582;
assign w584 = w559 & ~w583;
assign w585 = ~w559 & w583;
assign w586 = ~w584 & ~w585;
assign w587 = w532 & ~w586;
assign w588 = ~w532 & w586;
assign w589 = ~w587 & ~w588;
assign w590 = w520 & w589;
assign w591 = ~w520 & ~w589;
assign w592 = ~w590 & ~w591;
assign w593 = ~w518 & w592;
assign w594 = w518 & ~w592;
assign w595 = ~w593 & ~w594;
assign w596 = ~w503 & ~w595;
assign w597 = w503 & w595;
assign w598 = ~w596 & ~w597;
assign w599 = ~w507 & ~w510;
assign w600 = ~w513 & w8132;
assign w601 = (w598 & w513) | (w598 & w7499) | (w513 & w7499);
assign w602 = ~w600 & ~w601;
assign w603 = ~w530 & ~w586;
assign w604 = (~w527 & w529) | (~w527 & w7872) | (w529 & w7872);
assign w605 = ~w603 & w604;
assign w606 = w527 & w603;
assign w607 = ~w605 & ~w606;
assign w608 = (~w551 & ~w553) | (~w551 & w8133) | (~w553 & w8133);
assign w609 = w523 & w8134;
assign w610 = pi45 & w521;
assign w611 = ~pi45 & w522;
assign w612 = ~w610 & ~w611;
assign w613 = pi00 & ~w612;
assign w614 = pi01 & w523;
assign w615 = (w609 & w613) | (w609 & w8135) | (w613 & w8135);
assign w616 = ~w613 & w8136;
assign w617 = ~w615 & ~w616;
assign w618 = w608 & w617;
assign w619 = ~w608 & ~w617;
assign w620 = ~w618 & ~w619;
assign w621 = ~w558 & w583;
assign w622 = ~w557 & ~w621;
assign w623 = (w620 & w621) | (w620 & w8137) | (w621 & w8137);
assign w624 = ~w621 & w8138;
assign w625 = ~w623 & ~w624;
assign w626 = pi08 & ~w56;
assign w627 = pi09 & w56;
assign w628 = ~w626 & ~w627;
assign w629 = (~pi37 & w628) | (~pi37 & w7500) | (w628 & w7500);
assign w630 = w386 & ~w628;
assign w631 = ~w629 & ~w630;
assign w632 = pi10 & ~w25;
assign w633 = (pi35 & w632) | (pi35 & w7501) | (w632 & w7501);
assign w634 = ~w632 & w7502;
assign w635 = ~w633 & ~w634;
assign w636 = w631 & w635;
assign w637 = ~w631 & ~w635;
assign w638 = ~w636 & ~w637;
assign w639 = pi13 & pi32;
assign w640 = pi12 & ~pi32;
assign w641 = pi33 & ~w639;
assign w642 = ~w640 & w641;
assign w643 = ~pi33 & w639;
assign w644 = ~w642 & ~w643;
assign w645 = w638 & ~w644;
assign w646 = ~w638 & w644;
assign w647 = ~w645 & ~w646;
assign w648 = pi06 & ~w167;
assign w649 = pi07 & w119;
assign w650 = (pi39 & w648) | (pi39 & w8139) | (w648 & w8139);
assign w651 = ~w648 & w8140;
assign w652 = ~w650 & ~w651;
assign w653 = pi03 & w355;
assign w654 = (pi43 & ~w353) | (pi43 & w7503) | (~w353 & w7503);
assign w655 = w438 & w8141;
assign w656 = ~w653 & w8142;
assign w657 = pi43 & w653;
assign w658 = ~w656 & ~w657;
assign w659 = pi05 & w217;
assign w660 = (pi41 & ~w215) | (pi41 & w7504) | (~w215 & w7504);
assign w661 = w216 & w8143;
assign w662 = ~w659 & w8144;
assign w663 = pi41 & w659;
assign w664 = ~w662 & ~w663;
assign w665 = w658 & w664;
assign w666 = ~w658 & ~w664;
assign w667 = ~w665 & ~w666;
assign w668 = w652 & w667;
assign w669 = ~w652 & ~w667;
assign w670 = ~w668 & ~w669;
assign w671 = (~w572 & ~w574) | (~w572 & w7505) | (~w574 & w7505);
assign w672 = w670 & ~w671;
assign w673 = ~w670 & w671;
assign w674 = ~w672 & ~w673;
assign w675 = ~w647 & ~w674;
assign w676 = w647 & w674;
assign w677 = ~w675 & ~w676;
assign w678 = w625 & w677;
assign w679 = ~w625 & ~w677;
assign w680 = ~w678 & ~w679;
assign w681 = w607 & w680;
assign w682 = ~w607 & ~w680;
assign w683 = ~w681 & ~w682;
assign w684 = (w683 & w593) | (w683 & w8145) | (w593 & w8145);
assign w685 = ~w593 & w8146;
assign w686 = ~w684 & ~w685;
assign w687 = (w686 & w601) | (w686 & w8147) | (w601 & w8147);
assign w688 = ~w601 & w8148;
assign w689 = ~w687 & ~w688;
assign w690 = (pi45 & ~w523) | (pi45 & w8149) | (~w523 & w8149);
assign w691 = ~w613 & w8150;
assign w692 = ~w618 & ~w691;
assign w693 = ~w623 & ~w677;
assign w694 = ~w693 & w7506;
assign w695 = (w692 & w693) | (w692 & w7507) | (w693 & w7507);
assign w696 = ~w694 & ~w695;
assign w697 = (~w665 & ~w667) | (~w665 & w8151) | (~w667 & w8151);
assign w698 = ~pi45 & ~pi46;
assign w699 = pi45 & pi46;
assign w700 = ~w698 & ~w699;
assign w701 = pi00 & w700;
assign w702 = pi01 & ~w612;
assign w703 = (pi45 & w702) | (pi45 & w7873) | (w702 & w7873);
assign w704 = ~w702 & w7874;
assign w705 = ~w703 & ~w704;
assign w706 = w701 & w705;
assign w707 = ~w701 & ~w705;
assign w708 = ~w706 & ~w707;
assign w709 = ~w697 & w708;
assign w710 = w697 & ~w708;
assign w711 = ~w709 & ~w710;
assign w712 = (~w672 & ~w674) | (~w672 & w7508) | (~w674 & w7508);
assign w713 = w711 & ~w712;
assign w714 = ~w711 & w712;
assign w715 = ~w713 & ~w714;
assign w716 = pi07 & ~w167;
assign w717 = pi08 & w119;
assign w718 = (pi39 & w716) | (pi39 & w8152) | (w716 & w8152);
assign w719 = ~w716 & w8153;
assign w720 = ~w718 & ~w719;
assign w721 = pi05 & ~w304;
assign w722 = (pi41 & w721) | (pi41 & w7509) | (w721 & w7509);
assign w723 = ~w721 & w7510;
assign w724 = ~w722 & ~w723;
assign w725 = pi04 & w355;
assign w726 = (pi43 & ~w353) | (pi43 & w8154) | (~w353 & w8154);
assign w727 = pi03 & w354;
assign w728 = ~w725 & w8155;
assign w729 = pi43 & w725;
assign w730 = ~w728 & ~w729;
assign w731 = w724 & w730;
assign w732 = ~w724 & ~w730;
assign w733 = ~w731 & ~w732;
assign w734 = w720 & w733;
assign w735 = ~w720 & ~w733;
assign w736 = ~w734 & ~w735;
assign w737 = (~w636 & ~w638) | (~w636 & w7875) | (~w638 & w7875);
assign w738 = ~w736 & w737;
assign w739 = w736 & ~w737;
assign w740 = ~w738 & ~w739;
assign w741 = pi09 & ~w56;
assign w742 = pi10 & w56;
assign w743 = ~w741 & ~w742;
assign w744 = (~pi37 & w743) | (~pi37 & w7500) | (w743 & w7500);
assign w745 = w386 & ~w743;
assign w746 = ~w744 & ~w745;
assign w747 = pi11 & ~w25;
assign w748 = pi12 & w8;
assign w749 = (pi35 & w747) | (pi35 & w7511) | (w747 & w7511);
assign w750 = ~w747 & w7512;
assign w751 = ~w749 & ~w750;
assign w752 = w746 & w751;
assign w753 = ~w746 & ~w751;
assign w754 = ~w752 & ~w753;
assign w755 = pi14 & pi32;
assign w756 = pi13 & ~pi32;
assign w757 = pi33 & ~w755;
assign w758 = ~w756 & w757;
assign w759 = ~pi33 & w755;
assign w760 = ~w758 & ~w759;
assign w761 = w754 & ~w760;
assign w762 = ~w754 & w760;
assign w763 = ~w761 & ~w762;
assign w764 = w740 & ~w763;
assign w765 = ~w740 & w763;
assign w766 = ~w764 & ~w765;
assign w767 = w715 & ~w766;
assign w768 = ~w715 & w766;
assign w769 = ~w767 & ~w768;
assign w770 = w696 & ~w769;
assign w771 = ~w696 & w769;
assign w772 = ~w770 & ~w771;
assign w773 = (~w606 & ~w607) | (~w606 & w8156) | (~w607 & w8156);
assign w774 = ~w772 & ~w773;
assign w775 = w772 & w773;
assign w776 = ~w774 & ~w775;
assign w777 = (w601 & w8159) | (w601 & w8160) | (w8159 & w8160);
assign w778 = ~w776 & w9078;
assign w779 = ~w777 & ~w778;
assign w780 = ~w766 & w8161;
assign w781 = (~w709 & w712) | (~w709 & w7876) | (w712 & w7876);
assign w782 = (w781 & w766) | (w781 & w8162) | (w766 & w8162);
assign w783 = ~w780 & ~w782;
assign w784 = pi08 & ~w167;
assign w785 = pi09 & w119;
assign w786 = (pi39 & w784) | (pi39 & w8163) | (w784 & w8163);
assign w787 = ~w784 & w8164;
assign w788 = ~w786 & ~w787;
assign w789 = pi05 & w355;
assign w790 = ~pi42 & pi43;
assign w791 = ~w354 & ~w790;
assign w792 = pi41 & pi43;
assign w793 = pi04 & ~w792;
assign w794 = ~w791 & w793;
assign w795 = ~w789 & ~w794;
assign w796 = pi43 & ~w795;
assign w797 = ~pi43 & w795;
assign w798 = ~w796 & ~w797;
assign w799 = pi07 & w217;
assign w800 = ~pi40 & pi41;
assign w801 = ~w216 & ~w800;
assign w802 = pi39 & pi41;
assign w803 = pi06 & ~w802;
assign w804 = ~w801 & w803;
assign w805 = ~w799 & ~w804;
assign w806 = pi41 & ~w805;
assign w807 = ~pi41 & w805;
assign w808 = ~w806 & ~w807;
assign w809 = w798 & w808;
assign w810 = ~w798 & ~w808;
assign w811 = ~w809 & ~w810;
assign w812 = w788 & w811;
assign w813 = ~w788 & ~w811;
assign w814 = ~w812 & ~w813;
assign w815 = ~w753 & ~w760;
assign w816 = ~w752 & ~w815;
assign w817 = ~w814 & w816;
assign w818 = w814 & ~w816;
assign w819 = ~w817 & ~w818;
assign w820 = pi11 & w56;
assign w821 = (pi37 & ~w54) | (pi37 & w8165) | (~w54 & w8165);
assign w822 = pi10 & w55;
assign w823 = ~w820 & w8166;
assign w824 = pi37 & w820;
assign w825 = ~w823 & ~w824;
assign w826 = pi13 & w8;
assign w827 = (pi35 & ~w6) | (pi35 & w8167) | (~w6 & w8167);
assign w828 = pi12 & w7;
assign w829 = ~w826 & w8168;
assign w830 = pi35 & w826;
assign w831 = ~w829 & ~w830;
assign w832 = w825 & w831;
assign w833 = ~w825 & ~w831;
assign w834 = ~w832 & ~w833;
assign w835 = pi15 & pi32;
assign w836 = pi14 & ~pi32;
assign w837 = pi33 & ~w835;
assign w838 = ~w836 & w837;
assign w839 = ~pi33 & w835;
assign w840 = ~w838 & ~w839;
assign w841 = w834 & ~w840;
assign w842 = ~w834 & w840;
assign w843 = ~w841 & ~w842;
assign w844 = w819 & w843;
assign w845 = ~w819 & ~w843;
assign w846 = ~w844 & ~w845;
assign w847 = (~w731 & ~w733) | (~w731 & w8014) | (~w733 & w8014);
assign w848 = pi02 & ~w612;
assign w849 = (pi45 & w848) | (pi45 & w7513) | (w848 & w7513);
assign w850 = ~w848 & w7514;
assign w851 = ~w849 & ~w850;
assign w852 = ~pi47 & w699;
assign w853 = pi47 & w698;
assign w854 = ~w852 & ~w853;
assign w855 = pi00 & ~w854;
assign w856 = pi01 & w700;
assign w857 = (pi47 & w855) | (pi47 & w7515) | (w855 & w7515);
assign w858 = ~w855 & w7516;
assign w859 = ~w857 & ~w858;
assign w860 = w851 & w859;
assign w861 = ~w851 & ~w859;
assign w862 = ~w860 & ~w861;
assign w863 = (pi47 & ~w700) | (pi47 & w8169) | (~w700 & w8169);
assign w864 = (~w863 & ~w705) | (~w863 & w8015) | (~w705 & w8015);
assign w865 = w862 & ~w864;
assign w866 = ~w862 & w864;
assign w867 = ~w865 & ~w866;
assign w868 = ~w847 & w867;
assign w869 = w847 & ~w867;
assign w870 = ~w868 & ~w869;
assign w871 = ~w738 & w763;
assign w872 = ~w739 & ~w871;
assign w873 = w870 & ~w872;
assign w874 = ~w870 & w872;
assign w875 = ~w873 & ~w874;
assign w876 = w846 & ~w875;
assign w877 = ~w846 & w875;
assign w878 = ~w876 & ~w877;
assign w879 = w783 & ~w878;
assign w880 = ~w783 & w878;
assign w881 = ~w879 & ~w880;
assign w882 = ~w695 & ~w770;
assign w883 = ~w881 & ~w882;
assign w884 = w881 & w882;
assign w885 = ~w883 & ~w884;
assign w886 = ~w777 & w8170;
assign w887 = (~w885 & w777) | (~w885 & w8171) | (w777 & w8171);
assign w888 = ~w886 & ~w887;
assign w889 = ~w597 & ~w684;
assign w890 = ~w601 & w889;
assign w891 = w885 & w8172;
assign w892 = (~w780 & w878) | (~w780 & w8173) | (w878 & w8173);
assign w893 = (~w865 & ~w867) | (~w865 & w8016) | (~w867 & w8016);
assign w894 = ~pi49 & w893;
assign w895 = pi49 & ~w893;
assign w896 = ~w894 & ~w895;
assign w897 = w846 & ~w874;
assign w898 = (w896 & w897) | (w896 & w7877) | (w897 & w7877);
assign w899 = ~w897 & w7878;
assign w900 = ~w898 & ~w899;
assign w901 = (~w809 & ~w811) | (~w809 & w8174) | (~w811 & w8174);
assign w902 = pi03 & ~w612;
assign w903 = pi04 & w523;
assign w904 = (pi45 & w902) | (pi45 & w7517) | (w902 & w7517);
assign w905 = ~w902 & w7518;
assign w906 = ~w904 & ~w905;
assign w907 = ~pi47 & ~pi48;
assign w908 = pi47 & pi48;
assign w909 = ~w907 & ~w908;
assign w910 = (pi49 & ~w909) | (pi49 & w8175) | (~w909 & w8175);
assign w911 = w909 & w8176;
assign w912 = ~w910 & ~w911;
assign w913 = pi02 & w700;
assign w914 = (pi47 & ~w698) | (pi47 & w8177) | (~w698 & w8177);
assign w915 = pi01 & w699;
assign w916 = ~w913 & w8178;
assign w917 = pi47 & w913;
assign w918 = ~w916 & ~w917;
assign w919 = w912 & ~w918;
assign w920 = ~w912 & w918;
assign w921 = ~w919 & ~w920;
assign w922 = w860 & ~w921;
assign w923 = ~w860 & w921;
assign w924 = ~w922 & ~w923;
assign w925 = w906 & w924;
assign w926 = ~w906 & ~w924;
assign w927 = ~w925 & ~w926;
assign w928 = w901 & w927;
assign w929 = ~w901 & ~w927;
assign w930 = ~w928 & ~w929;
assign w931 = (~w818 & ~w819) | (~w818 & w7519) | (~w819 & w7519);
assign w932 = w930 & ~w931;
assign w933 = ~w930 & w931;
assign w934 = ~w932 & ~w933;
assign w935 = (~w832 & ~w834) | (~w832 & w7520) | (~w834 & w7520);
assign w936 = pi09 & ~w167;
assign w937 = pi10 & w119;
assign w938 = (pi39 & w936) | (pi39 & w7521) | (w936 & w7521);
assign w939 = ~w936 & w7522;
assign w940 = ~w938 & ~w939;
assign w941 = pi08 & w217;
assign w942 = (pi41 & ~w215) | (pi41 & w8179) | (~w215 & w8179);
assign w943 = pi07 & w216;
assign w944 = ~w941 & w8180;
assign w945 = pi41 & w941;
assign w946 = ~w944 & ~w945;
assign w947 = pi06 & w355;
assign w948 = (pi43 & ~w353) | (pi43 & w8181) | (~w353 & w8181);
assign w949 = pi05 & w354;
assign w950 = ~w947 & w8182;
assign w951 = pi43 & w947;
assign w952 = ~w950 & ~w951;
assign w953 = ~w946 & ~w952;
assign w954 = w946 & w952;
assign w955 = ~w953 & ~w954;
assign w956 = w940 & w955;
assign w957 = ~w940 & ~w955;
assign w958 = ~w956 & ~w957;
assign w959 = ~w935 & w958;
assign w960 = w935 & ~w958;
assign w961 = ~w959 & ~w960;
assign w962 = pi14 & w8;
assign w963 = (pi35 & ~w6) | (pi35 & w8183) | (~w6 & w8183);
assign w964 = pi13 & w7;
assign w965 = ~w962 & w8184;
assign w966 = pi35 & w962;
assign w967 = ~w965 & ~w966;
assign w968 = pi12 & w56;
assign w969 = (pi37 & ~w54) | (pi37 & w8185) | (~w54 & w8185);
assign w970 = pi11 & w55;
assign w971 = ~w968 & w8186;
assign w972 = pi37 & w968;
assign w973 = ~w971 & ~w972;
assign w974 = w967 & w973;
assign w975 = ~w967 & ~w973;
assign w976 = ~w974 & ~w975;
assign w977 = pi16 & pi32;
assign w978 = pi15 & ~pi32;
assign w979 = pi33 & ~w977;
assign w980 = ~w978 & w979;
assign w981 = ~pi33 & w977;
assign w982 = ~w980 & ~w981;
assign w983 = w976 & ~w982;
assign w984 = ~w976 & w982;
assign w985 = ~w983 & ~w984;
assign w986 = w961 & w985;
assign w987 = ~w961 & ~w985;
assign w988 = ~w986 & ~w987;
assign w989 = w934 & w988;
assign w990 = ~w934 & ~w988;
assign w991 = ~w989 & ~w990;
assign w992 = ~w900 & ~w991;
assign w993 = w900 & w991;
assign w994 = ~w992 & ~w993;
assign w995 = w892 & ~w994;
assign w996 = ~w892 & w994;
assign w997 = ~w995 & ~w996;
assign w998 = ~w774 & ~w884;
assign w999 = ~w883 & ~w998;
assign w1000 = w997 & w999;
assign w1001 = ~w997 & ~w999;
assign w1002 = ~w1000 & ~w1001;
assign w1003 = (~w1002 & w890) | (~w1002 & w8187) | (w890 & w8187);
assign w1004 = ~w890 & w1122;
assign w1005 = ~w1003 & ~w1004;
assign w1006 = ~w884 & ~w996;
assign w1007 = ~w995 & ~w1006;
assign w1008 = w860 & w927;
assign w1009 = ~w929 & ~w1008;
assign w1010 = ~w932 & ~w988;
assign w1011 = (w1009 & w1010) | (w1009 & w7523) | (w1010 & w7523);
assign w1012 = ~w1010 & w7524;
assign w1013 = ~w1011 & ~w1012;
assign w1014 = ~w940 & ~w954;
assign w1015 = ~w953 & ~w1014;
assign w1016 = ~w906 & ~w920;
assign w1017 = ~w919 & ~w1016;
assign w1018 = w1015 & w1017;
assign w1019 = ~w1015 & ~w1017;
assign w1020 = ~w1018 & ~w1019;
assign w1021 = pi04 & ~w612;
assign w1022 = (pi45 & w1021) | (pi45 & w7525) | (w1021 & w7525);
assign w1023 = ~w1021 & w7526;
assign w1024 = ~w1022 & ~w1023;
assign w1025 = pi03 & w700;
assign w1026 = (pi47 & ~w698) | (pi47 & w8188) | (~w698 & w8188);
assign w1027 = pi02 & w699;
assign w1028 = ~w1025 & w8189;
assign w1029 = w700 & w8998;
assign w1030 = ~w1028 & ~w1029;
assign w1031 = pi01 & w909;
assign w1032 = (pi49 & ~w907) | (pi49 & w8175) | (~w907 & w8175);
assign w1033 = pi00 & w908;
assign w1034 = ~w1031 & w8190;
assign w1035 = w909 & w8999;
assign w1036 = ~w1034 & ~w1035;
assign w1037 = w1030 & w1036;
assign w1038 = ~w1030 & ~w1036;
assign w1039 = ~w1037 & ~w1038;
assign w1040 = w1024 & w1039;
assign w1041 = ~w1024 & ~w1039;
assign w1042 = ~w1040 & ~w1041;
assign w1043 = w1020 & w1042;
assign w1044 = ~w1020 & ~w1042;
assign w1045 = ~w1043 & ~w1044;
assign w1046 = ~w959 & ~w985;
assign w1047 = ~w960 & ~w1046;
assign w1048 = w1045 & w1047;
assign w1049 = ~w1045 & ~w1047;
assign w1050 = ~w1048 & ~w1049;
assign w1051 = (~w974 & ~w976) | (~w974 & w7527) | (~w976 & w7527);
assign w1052 = pi10 & ~w167;
assign w1053 = (pi39 & w1052) | (pi39 & w7528) | (w1052 & w7528);
assign w1054 = ~w1052 & w7529;
assign w1055 = ~w1053 & ~w1054;
assign w1056 = pi09 & w217;
assign w1057 = (pi41 & ~w215) | (pi41 & w8191) | (~w215 & w8191);
assign w1058 = pi08 & w216;
assign w1059 = ~w1056 & w8192;
assign w1060 = w217 & w9000;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = pi07 & w355;
assign w1063 = (pi43 & ~w353) | (pi43 & w8193) | (~w353 & w8193);
assign w1064 = pi06 & w354;
assign w1065 = ~w1062 & w8194;
assign w1066 = w355 & w9001;
assign w1067 = ~w1065 & ~w1066;
assign w1068 = ~w1061 & ~w1067;
assign w1069 = w1061 & w1067;
assign w1070 = ~w1068 & ~w1069;
assign w1071 = w1055 & w1070;
assign w1072 = ~w1055 & ~w1070;
assign w1073 = ~w1071 & ~w1072;
assign w1074 = ~w1051 & w1073;
assign w1075 = w1051 & ~w1073;
assign w1076 = ~w1074 & ~w1075;
assign w1077 = pi13 & w56;
assign w1078 = (pi37 & ~w54) | (pi37 & w8195) | (~w54 & w8195);
assign w1079 = pi12 & w55;
assign w1080 = ~w1077 & w8196;
assign w1081 = pi37 & w1077;
assign w1082 = ~w1080 & ~w1081;
assign w1083 = pi15 & w8;
assign w1084 = (pi35 & ~w6) | (pi35 & w8197) | (~w6 & w8197);
assign w1085 = pi14 & w7;
assign w1086 = ~w1083 & w8198;
assign w1087 = pi35 & w1083;
assign w1088 = ~w1086 & ~w1087;
assign w1089 = w1082 & w1088;
assign w1090 = ~w1082 & ~w1088;
assign w1091 = ~w1089 & ~w1090;
assign w1092 = pi17 & pi32;
assign w1093 = pi16 & ~pi32;
assign w1094 = pi33 & ~w1092;
assign w1095 = ~w1093 & w1094;
assign w1096 = ~pi33 & w1092;
assign w1097 = ~w1095 & ~w1096;
assign w1098 = w1091 & ~w1097;
assign w1099 = ~w1091 & w1097;
assign w1100 = ~w1098 & ~w1099;
assign w1101 = w1076 & w1100;
assign w1102 = ~w1076 & ~w1100;
assign w1103 = ~w1101 & ~w1102;
assign w1104 = w1050 & w1103;
assign w1105 = ~w1050 & ~w1103;
assign w1106 = ~w1104 & ~w1105;
assign w1107 = w1013 & w1106;
assign w1108 = ~w1013 & ~w1106;
assign w1109 = ~w1107 & ~w1108;
assign w1110 = w991 & w7879;
assign w1111 = ~w895 & ~w898;
assign w1112 = (w1111 & ~w991) | (w1111 & w7880) | (~w991 & w7880);
assign w1113 = ~w1110 & ~w1112;
assign w1114 = w1109 & w1113;
assign w1115 = ~w1109 & ~w1113;
assign w1116 = ~w1114 & ~w1115;
assign w1117 = w1007 & w1116;
assign w1118 = ~w1007 & ~w1116;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = w999 & w8199;
assign w1121 = w1119 & w1120;
assign w1122 = w891 & w1002;
assign w1123 = w1119 & w1122;
assign w1124 = ~w890 & w1123;
assign w1125 = ~w1119 & ~w1120;
assign w1126 = ~w1004 & w1125;
assign w1127 = (~w1121 & ~w1123) | (~w1121 & w8200) | (~w1123 & w8200);
assign w1128 = ~w1126 & w1127;
assign w1129 = (~w1012 & ~w1013) | (~w1012 & w8017) | (~w1013 & w8017);
assign w1130 = ~pi49 & ~pi50;
assign w1131 = pi49 & pi50;
assign w1132 = ~w1130 & ~w1131;
assign w1133 = pi00 & w1132;
assign w1134 = (~w1018 & ~w1020) | (~w1018 & w8201) | (~w1020 & w8201);
assign w1135 = w1133 & ~w1134;
assign w1136 = ~w1133 & w1134;
assign w1137 = ~w1135 & ~w1136;
assign w1138 = ~w1048 & ~w1103;
assign w1139 = ~w1049 & ~w1138;
assign w1140 = (~w1137 & w1138) | (~w1137 & w8202) | (w1138 & w8202);
assign w1141 = ~w1138 & w8203;
assign w1142 = ~w1140 & ~w1141;
assign w1143 = ~w1024 & ~w1037;
assign w1144 = ~w1038 & ~w1143;
assign w1145 = ~w1055 & ~w1069;
assign w1146 = ~w1068 & ~w1145;
assign w1147 = w1144 & w1146;
assign w1148 = ~w1144 & ~w1146;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = pi05 & ~w612;
assign w1151 = (pi45 & w1150) | (pi45 & w7530) | (w1150 & w7530);
assign w1152 = ~w1150 & w7531;
assign w1153 = ~w1151 & ~w1152;
assign w1154 = pi04 & w700;
assign w1155 = (pi47 & ~w698) | (pi47 & w8204) | (~w698 & w8204);
assign w1156 = pi03 & w699;
assign w1157 = ~w1154 & w8205;
assign w1158 = w700 & w9002;
assign w1159 = ~w1157 & ~w1158;
assign w1160 = pi02 & w909;
assign w1161 = (pi49 & ~w907) | (pi49 & w8206) | (~w907 & w8206);
assign w1162 = pi01 & w908;
assign w1163 = ~w1160 & w8207;
assign w1164 = w909 & w9003;
assign w1165 = ~w1163 & ~w1164;
assign w1166 = w1159 & w1165;
assign w1167 = ~w1159 & ~w1165;
assign w1168 = ~w1166 & ~w1167;
assign w1169 = w1153 & w1168;
assign w1170 = ~w1153 & ~w1168;
assign w1171 = ~w1169 & ~w1170;
assign w1172 = ~w1149 & ~w1171;
assign w1173 = w1149 & w1171;
assign w1174 = ~w1172 & ~w1173;
assign w1175 = ~w1074 & ~w1100;
assign w1176 = ~w1075 & ~w1175;
assign w1177 = w1174 & w1176;
assign w1178 = ~w1174 & ~w1176;
assign w1179 = ~w1177 & ~w1178;
assign w1180 = (~w1089 & ~w1091) | (~w1089 & w7532) | (~w1091 & w7532);
assign w1181 = pi11 & ~w167;
assign w1182 = (pi39 & w1181) | (pi39 & w7533) | (w1181 & w7533);
assign w1183 = ~w1181 & w7534;
assign w1184 = ~w1182 & ~w1183;
assign w1185 = pi10 & w217;
assign w1186 = (pi41 & ~w215) | (pi41 & w8208) | (~w215 & w8208);
assign w1187 = pi09 & w216;
assign w1188 = ~w1185 & w8209;
assign w1189 = w217 & w9004;
assign w1190 = ~w1188 & ~w1189;
assign w1191 = pi08 & w355;
assign w1192 = (pi43 & ~w353) | (pi43 & w8210) | (~w353 & w8210);
assign w1193 = pi07 & w354;
assign w1194 = ~w1191 & w8211;
assign w1195 = w355 & w9005;
assign w1196 = ~w1194 & ~w1195;
assign w1197 = ~w1190 & ~w1196;
assign w1198 = w1190 & w1196;
assign w1199 = ~w1197 & ~w1198;
assign w1200 = w1184 & w1199;
assign w1201 = ~w1184 & ~w1199;
assign w1202 = ~w1200 & ~w1201;
assign w1203 = ~w1180 & w1202;
assign w1204 = w1180 & ~w1202;
assign w1205 = ~w1203 & ~w1204;
assign w1206 = pi16 & w8;
assign w1207 = (pi35 & ~w6) | (pi35 & w8212) | (~w6 & w8212);
assign w1208 = pi15 & w7;
assign w1209 = ~w1206 & w8213;
assign w1210 = pi35 & w1206;
assign w1211 = ~w1209 & ~w1210;
assign w1212 = pi14 & w56;
assign w1213 = (pi37 & ~w54) | (pi37 & w8214) | (~w54 & w8214);
assign w1214 = pi13 & w55;
assign w1215 = ~w1212 & w8215;
assign w1216 = pi37 & w1212;
assign w1217 = ~w1215 & ~w1216;
assign w1218 = w1211 & w1217;
assign w1219 = ~w1211 & ~w1217;
assign w1220 = ~w1218 & ~w1219;
assign w1221 = pi18 & pi32;
assign w1222 = pi17 & ~pi32;
assign w1223 = pi33 & ~w1221;
assign w1224 = ~w1222 & w1223;
assign w1225 = ~pi33 & w1221;
assign w1226 = ~w1224 & ~w1225;
assign w1227 = w1220 & ~w1226;
assign w1228 = ~w1220 & w1226;
assign w1229 = ~w1227 & ~w1228;
assign w1230 = w1205 & w1229;
assign w1231 = ~w1205 & ~w1229;
assign w1232 = ~w1230 & ~w1231;
assign w1233 = w1179 & w1232;
assign w1234 = ~w1179 & ~w1232;
assign w1235 = ~w1233 & ~w1234;
assign w1236 = w1142 & ~w1235;
assign w1237 = ~w1142 & w1235;
assign w1238 = ~w1236 & ~w1237;
assign w1239 = ~w1129 & ~w1238;
assign w1240 = w1129 & w1238;
assign w1241 = ~w1239 & ~w1240;
assign w1242 = (~w1110 & ~w1113) | (~w1110 & w8216) | (~w1113 & w8216);
assign w1243 = w1241 & ~w1242;
assign w1244 = ~w1241 & w1242;
assign w1245 = ~w1243 & ~w1244;
assign w1246 = (~w1117 & ~w1119) | (~w1117 & w7881) | (~w1119 & w7881);
assign w1247 = (w1246 & ~w1123) | (w1246 & w8217) | (~w1123 & w8217);
assign w1248 = ~w1245 & w1247;
assign w1249 = w1245 & ~w1247;
assign w1250 = ~w1248 & ~w1249;
assign w1251 = ~w1140 & w1235;
assign w1252 = (~w1135 & ~w1139) | (~w1135 & w7535) | (~w1139 & w7535);
assign w1253 = ~w1251 & w1252;
assign w1254 = w1235 & w8218;
assign w1255 = ~w1253 & ~w1254;
assign w1256 = (~w1147 & ~w1149) | (~w1147 & w8219) | (~w1149 & w8219);
assign w1257 = w1132 & w8220;
assign w1258 = pi51 & w1130;
assign w1259 = ~pi51 & w1131;
assign w1260 = ~w1258 & ~w1259;
assign w1261 = pi00 & ~w1260;
assign w1262 = pi01 & w1132;
assign w1263 = (w1257 & w1261) | (w1257 & w8221) | (w1261 & w8221);
assign w1264 = ~w1261 & w8222;
assign w1265 = ~w1263 & ~w1264;
assign w1266 = ~w1256 & w1265;
assign w1267 = w1256 & ~w1265;
assign w1268 = ~w1266 & ~w1267;
assign w1269 = ~w1177 & ~w1232;
assign w1270 = ~w1178 & ~w1269;
assign w1271 = (~w1268 & w1269) | (~w1268 & w8223) | (w1269 & w8223);
assign w1272 = ~w1269 & w8224;
assign w1273 = ~w1271 & ~w1272;
assign w1274 = ~w1153 & ~w1166;
assign w1275 = ~w1167 & ~w1274;
assign w1276 = ~w1184 & ~w1198;
assign w1277 = ~w1197 & ~w1276;
assign w1278 = w1275 & w1277;
assign w1279 = ~w1275 & ~w1277;
assign w1280 = ~w1278 & ~w1279;
assign w1281 = pi06 & ~w612;
assign w1282 = pi07 & w523;
assign w1283 = (pi45 & w1281) | (pi45 & w7536) | (w1281 & w7536);
assign w1284 = ~w1281 & w7537;
assign w1285 = ~w1283 & ~w1284;
assign w1286 = pi05 & w700;
assign w1287 = (pi47 & ~w698) | (pi47 & w8225) | (~w698 & w8225);
assign w1288 = pi04 & w699;
assign w1289 = ~w1286 & w8226;
assign w1290 = pi47 & w1286;
assign w1291 = ~w1289 & ~w1290;
assign w1292 = pi03 & w909;
assign w1293 = (pi49 & ~w907) | (pi49 & w8227) | (~w907 & w8227);
assign w1294 = pi02 & w908;
assign w1295 = ~w1292 & w8228;
assign w1296 = pi49 & w1292;
assign w1297 = ~w1295 & ~w1296;
assign w1298 = w1291 & w1297;
assign w1299 = ~w1291 & ~w1297;
assign w1300 = ~w1298 & ~w1299;
assign w1301 = w1285 & w1300;
assign w1302 = ~w1285 & ~w1300;
assign w1303 = ~w1301 & ~w1302;
assign w1304 = w1280 & ~w1303;
assign w1305 = ~w1280 & w1303;
assign w1306 = ~w1304 & ~w1305;
assign w1307 = ~w1203 & ~w1229;
assign w1308 = ~w1204 & ~w1307;
assign w1309 = w1306 & ~w1308;
assign w1310 = ~w1306 & w1308;
assign w1311 = ~w1309 & ~w1310;
assign w1312 = (~w1218 & ~w1220) | (~w1218 & w7538) | (~w1220 & w7538);
assign w1313 = pi12 & ~w167;
assign w1314 = pi13 & w119;
assign w1315 = (pi39 & w1313) | (pi39 & w7539) | (w1313 & w7539);
assign w1316 = ~w1313 & w7540;
assign w1317 = ~w1315 & ~w1316;
assign w1318 = pi11 & w217;
assign w1319 = (pi41 & ~w215) | (pi41 & w8229) | (~w215 & w8229);
assign w1320 = pi10 & w216;
assign w1321 = ~w1318 & w8230;
assign w1322 = pi41 & w1318;
assign w1323 = ~w1321 & ~w1322;
assign w1324 = pi09 & w355;
assign w1325 = (pi43 & ~w353) | (pi43 & w8231) | (~w353 & w8231);
assign w1326 = pi08 & w354;
assign w1327 = ~w1324 & w8232;
assign w1328 = pi43 & w1324;
assign w1329 = ~w1327 & ~w1328;
assign w1330 = ~w1323 & ~w1329;
assign w1331 = w1323 & w1329;
assign w1332 = ~w1330 & ~w1331;
assign w1333 = w1317 & w1332;
assign w1334 = ~w1317 & ~w1332;
assign w1335 = ~w1333 & ~w1334;
assign w1336 = ~w1312 & w1335;
assign w1337 = w1312 & ~w1335;
assign w1338 = ~w1336 & ~w1337;
assign w1339 = pi15 & w56;
assign w1340 = (pi37 & ~w54) | (pi37 & w8233) | (~w54 & w8233);
assign w1341 = pi14 & w55;
assign w1342 = ~w1339 & w8234;
assign w1343 = pi37 & w1339;
assign w1344 = ~w1342 & ~w1343;
assign w1345 = pi17 & w8;
assign w1346 = (pi35 & ~w6) | (pi35 & w8235) | (~w6 & w8235);
assign w1347 = pi16 & w7;
assign w1348 = ~w1345 & w8236;
assign w1349 = pi35 & w1345;
assign w1350 = ~w1348 & ~w1349;
assign w1351 = w1344 & w1350;
assign w1352 = ~w1344 & ~w1350;
assign w1353 = ~w1351 & ~w1352;
assign w1354 = pi19 & pi32;
assign w1355 = pi18 & ~pi32;
assign w1356 = pi33 & ~w1354;
assign w1357 = ~w1355 & w1356;
assign w1358 = ~pi33 & w1354;
assign w1359 = ~w1357 & ~w1358;
assign w1360 = w1353 & ~w1359;
assign w1361 = ~w1353 & w1359;
assign w1362 = ~w1360 & ~w1361;
assign w1363 = w1338 & w1362;
assign w1364 = ~w1338 & ~w1362;
assign w1365 = ~w1363 & ~w1364;
assign w1366 = w1311 & w1365;
assign w1367 = ~w1311 & ~w1365;
assign w1368 = ~w1366 & ~w1367;
assign w1369 = w1273 & ~w1368;
assign w1370 = ~w1273 & w1368;
assign w1371 = ~w1369 & ~w1370;
assign w1372 = w1255 & w1371;
assign w1373 = ~w1255 & ~w1371;
assign w1374 = ~w1372 & ~w1373;
assign w1375 = ~w1239 & w1374;
assign w1376 = w1239 & ~w1374;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = ~w1243 & ~w1377;
assign w1379 = w1243 & ~w1374;
assign w1380 = w1245 & w1377;
assign w1381 = (~w1379 & w1247) | (~w1379 & w8237) | (w1247 & w8237);
assign w1382 = ~w1378 & w1381;
assign w1383 = ~w1247 & w8238;
assign w1384 = ~w1382 & ~w1383;
assign w1385 = (~w1253 & ~w1255) | (~w1253 & w8239) | (~w1255 & w8239);
assign w1386 = ~w1271 & w1368;
assign w1387 = w1368 & w8240;
assign w1388 = (~w1266 & ~w1270) | (~w1266 & w7541) | (~w1270 & w7541);
assign w1389 = ~w1386 & w1388;
assign w1390 = ~w1387 & ~w1389;
assign w1391 = ~pi51 & ~pi52;
assign w1392 = pi51 & pi52;
assign w1393 = ~w1391 & ~w1392;
assign w1394 = pi00 & w1393;
assign w1395 = pi02 & w1132;
assign w1396 = (pi51 & ~w1130) | (pi51 & w8241) | (~w1130 & w8241);
assign w1397 = pi01 & w1131;
assign w1398 = ~w1395 & w8242;
assign w1399 = pi51 & w1395;
assign w1400 = ~w1398 & ~w1399;
assign w1401 = w1394 & ~w1400;
assign w1402 = ~w1394 & w1400;
assign w1403 = ~w1401 & ~w1402;
assign w1404 = (pi51 & ~w1132) | (pi51 & w8243) | (~w1132 & w8243);
assign w1405 = ~w1261 & w8244;
assign w1406 = w1403 & ~w1405;
assign w1407 = ~w1403 & w1405;
assign w1408 = ~w1406 & ~w1407;
assign w1409 = (~w1279 & ~w1280) | (~w1279 & w8245) | (~w1280 & w8245);
assign w1410 = w1408 & w1409;
assign w1411 = ~w1408 & ~w1409;
assign w1412 = ~w1410 & ~w1411;
assign w1413 = ~w1310 & ~w1365;
assign w1414 = ~w1309 & ~w1413;
assign w1415 = ~w1413 & w8246;
assign w1416 = (~w1412 & w1413) | (~w1412 & w8247) | (w1413 & w8247);
assign w1417 = ~w1415 & ~w1416;
assign w1418 = ~w1285 & ~w1298;
assign w1419 = ~w1299 & ~w1418;
assign w1420 = ~w1317 & ~w1331;
assign w1421 = ~w1330 & ~w1420;
assign w1422 = w1419 & w1421;
assign w1423 = ~w1419 & ~w1421;
assign w1424 = ~w1422 & ~w1423;
assign w1425 = pi07 & ~w612;
assign w1426 = (pi45 & w1425) | (pi45 & w7542) | (w1425 & w7542);
assign w1427 = ~w1425 & w7543;
assign w1428 = ~w1426 & ~w1427;
assign w1429 = pi06 & w700;
assign w1430 = (pi47 & ~w698) | (pi47 & w8248) | (~w698 & w8248);
assign w1431 = pi05 & w699;
assign w1432 = ~w1429 & w8249;
assign w1433 = w700 & w9006;
assign w1434 = ~w1432 & ~w1433;
assign w1435 = pi04 & w909;
assign w1436 = (pi49 & ~w907) | (pi49 & w8250) | (~w907 & w8250);
assign w1437 = pi03 & w908;
assign w1438 = ~w1435 & w8251;
assign w1439 = w909 & w9007;
assign w1440 = ~w1438 & ~w1439;
assign w1441 = w1434 & w1440;
assign w1442 = ~w1434 & ~w1440;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = w1428 & w1443;
assign w1445 = ~w1428 & ~w1443;
assign w1446 = ~w1444 & ~w1445;
assign w1447 = ~w1424 & ~w1446;
assign w1448 = w1424 & w1446;
assign w1449 = ~w1447 & ~w1448;
assign w1450 = ~w1336 & ~w1362;
assign w1451 = ~w1337 & ~w1450;
assign w1452 = w1449 & w1451;
assign w1453 = ~w1449 & ~w1451;
assign w1454 = ~w1452 & ~w1453;
assign w1455 = (~w1351 & ~w1353) | (~w1351 & w7544) | (~w1353 & w7544);
assign w1456 = pi13 & ~w167;
assign w1457 = (pi39 & w1456) | (pi39 & w7545) | (w1456 & w7545);
assign w1458 = ~w1456 & w7546;
assign w1459 = ~w1457 & ~w1458;
assign w1460 = pi12 & w217;
assign w1461 = (pi41 & ~w215) | (pi41 & w8252) | (~w215 & w8252);
assign w1462 = pi11 & w216;
assign w1463 = ~w1460 & w8253;
assign w1464 = w217 & w9008;
assign w1465 = ~w1463 & ~w1464;
assign w1466 = pi10 & w355;
assign w1467 = (pi43 & ~w353) | (pi43 & w8254) | (~w353 & w8254);
assign w1468 = pi09 & w354;
assign w1469 = ~w1466 & w8255;
assign w1470 = w355 & w9009;
assign w1471 = ~w1469 & ~w1470;
assign w1472 = ~w1465 & ~w1471;
assign w1473 = w1465 & w1471;
assign w1474 = ~w1472 & ~w1473;
assign w1475 = w1459 & w1474;
assign w1476 = ~w1459 & ~w1474;
assign w1477 = ~w1475 & ~w1476;
assign w1478 = ~w1455 & w1477;
assign w1479 = w1455 & ~w1477;
assign w1480 = ~w1478 & ~w1479;
assign w1481 = pi18 & w8;
assign w1482 = (pi35 & ~w6) | (pi35 & w8256) | (~w6 & w8256);
assign w1483 = pi17 & w7;
assign w1484 = ~w1481 & w8257;
assign w1485 = pi35 & w1481;
assign w1486 = ~w1484 & ~w1485;
assign w1487 = pi16 & w56;
assign w1488 = (pi37 & ~w54) | (pi37 & w8258) | (~w54 & w8258);
assign w1489 = pi15 & w55;
assign w1490 = ~w1487 & w8259;
assign w1491 = pi37 & w1487;
assign w1492 = ~w1490 & ~w1491;
assign w1493 = w1486 & w1492;
assign w1494 = ~w1486 & ~w1492;
assign w1495 = ~w1493 & ~w1494;
assign w1496 = pi20 & pi32;
assign w1497 = pi19 & ~pi32;
assign w1498 = pi33 & ~w1496;
assign w1499 = ~w1497 & w1498;
assign w1500 = ~pi33 & w1496;
assign w1501 = ~w1499 & ~w1500;
assign w1502 = w1495 & ~w1501;
assign w1503 = ~w1495 & w1501;
assign w1504 = ~w1502 & ~w1503;
assign w1505 = w1480 & w1504;
assign w1506 = ~w1480 & ~w1504;
assign w1507 = ~w1505 & ~w1506;
assign w1508 = w1454 & ~w1507;
assign w1509 = ~w1454 & w1507;
assign w1510 = ~w1508 & ~w1509;
assign w1511 = w1417 & ~w1510;
assign w1512 = ~w1417 & w1510;
assign w1513 = ~w1511 & ~w1512;
assign w1514 = w1390 & w1513;
assign w1515 = ~w1390 & ~w1513;
assign w1516 = ~w1514 & ~w1515;
assign w1517 = w1385 & w1516;
assign w1518 = ~w1385 & ~w1516;
assign w1519 = ~w1517 & ~w1518;
assign w1520 = w1380 & w1519;
assign w1521 = ~w1376 & ~w1519;
assign w1522 = w1376 & w1519;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = w1379 & w1523;
assign w1525 = ~w1524 & w9092;
assign w1526 = w1381 & ~w1523;
assign w1527 = w1525 & ~w1526;
assign w1528 = (~w1387 & ~w1390) | (~w1387 & w8260) | (~w1390 & w8260);
assign w1529 = (~w1407 & ~w1409) | (~w1407 & w8261) | (~w1409 & w8261);
assign w1530 = ~w1415 & w1510;
assign w1531 = (w1529 & w1530) | (w1529 & w7547) | (w1530 & w7547);
assign w1532 = ~w1530 & w7548;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = ~pi53 & w1392;
assign w1535 = pi53 & w1391;
assign w1536 = ~w1534 & ~w1535;
assign w1537 = pi00 & ~w1536;
assign w1538 = pi01 & w1393;
assign w1539 = (pi53 & w1537) | (pi53 & w7549) | (w1537 & w7549);
assign w1540 = ~w1537 & w7550;
assign w1541 = ~w1539 & ~w1540;
assign w1542 = pi02 & ~w1260;
assign w1543 = pi03 & w1132;
assign w1544 = (pi51 & w1542) | (pi51 & w7551) | (w1542 & w7551);
assign w1545 = ~w1542 & w7552;
assign w1546 = ~w1544 & ~w1545;
assign w1547 = w1541 & w1546;
assign w1548 = ~w1541 & ~w1546;
assign w1549 = ~w1547 & ~w1548;
assign w1550 = (~pi53 & ~w1393) | (~pi53 & w8262) | (~w1393 & w8262);
assign w1551 = (~w1550 & w1400) | (~w1550 & w8263) | (w1400 & w8263);
assign w1552 = ~w1549 & ~w1551;
assign w1553 = w1549 & w1551;
assign w1554 = ~w1552 & ~w1553;
assign w1555 = (~w1422 & ~w1424) | (~w1422 & w8264) | (~w1424 & w8264);
assign w1556 = w1554 & ~w1555;
assign w1557 = ~w1554 & w1555;
assign w1558 = ~w1556 & ~w1557;
assign w1559 = (~w1453 & ~w1454) | (~w1453 & w7553) | (~w1454 & w7553);
assign w1560 = ~w1428 & ~w1441;
assign w1561 = ~w1442 & ~w1560;
assign w1562 = ~w1459 & ~w1473;
assign w1563 = ~w1472 & ~w1562;
assign w1564 = w1561 & w1563;
assign w1565 = ~w1561 & ~w1563;
assign w1566 = ~w1564 & ~w1565;
assign w1567 = pi09 & w523;
assign w1568 = ~pi44 & pi45;
assign w1569 = ~w522 & ~w1568;
assign w1570 = pi43 & pi45;
assign w1571 = pi08 & ~w1570;
assign w1572 = ~w1569 & w1571;
assign w1573 = ~w1567 & ~w1572;
assign w1574 = pi45 & ~w1573;
assign w1575 = ~pi45 & w1573;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = pi07 & w700;
assign w1578 = (pi47 & ~w698) | (pi47 & w8265) | (~w698 & w8265);
assign w1579 = pi06 & w699;
assign w1580 = ~w1577 & w8266;
assign w1581 = pi47 & w1577;
assign w1582 = ~w1580 & ~w1581;
assign w1583 = ~w1576 & ~w1582;
assign w1584 = w1576 & w1582;
assign w1585 = ~w1583 & ~w1584;
assign w1586 = pi05 & w909;
assign w1587 = (pi49 & ~w907) | (pi49 & w8267) | (~w907 & w8267);
assign w1588 = pi04 & w908;
assign w1589 = ~w1586 & w8268;
assign w1590 = pi49 & w1586;
assign w1591 = ~w1589 & ~w1590;
assign w1592 = w1585 & ~w1591;
assign w1593 = ~w1585 & w1591;
assign w1594 = ~w1592 & ~w1593;
assign w1595 = ~w1566 & w1594;
assign w1596 = w1566 & ~w1594;
assign w1597 = ~w1595 & ~w1596;
assign w1598 = ~w1478 & ~w1504;
assign w1599 = ~w1479 & ~w1598;
assign w1600 = w1597 & w1599;
assign w1601 = ~w1597 & ~w1599;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = (~w1493 & ~w1495) | (~w1493 & w7554) | (~w1495 & w7554);
assign w1604 = pi19 & w8;
assign w1605 = (pi35 & ~w6) | (pi35 & w8269) | (~w6 & w8269);
assign w1606 = pi18 & w7;
assign w1607 = ~w1604 & w8270;
assign w1608 = pi35 & w1604;
assign w1609 = ~w1607 & ~w1608;
assign w1610 = pi17 & w56;
assign w1611 = (pi37 & ~w54) | (pi37 & w8271) | (~w54 & w8271);
assign w1612 = pi16 & w55;
assign w1613 = ~w1610 & w8272;
assign w1614 = pi37 & w1610;
assign w1615 = ~w1613 & ~w1614;
assign w1616 = w1609 & w1615;
assign w1617 = ~w1609 & ~w1615;
assign w1618 = ~w1616 & ~w1617;
assign w1619 = pi21 & pi32;
assign w1620 = pi20 & ~pi32;
assign w1621 = pi33 & ~w1619;
assign w1622 = ~w1620 & w1621;
assign w1623 = ~pi33 & w1619;
assign w1624 = ~w1622 & ~w1623;
assign w1625 = w1618 & ~w1624;
assign w1626 = ~w1618 & w1624;
assign w1627 = ~w1625 & ~w1626;
assign w1628 = ~w1603 & w1627;
assign w1629 = w1603 & ~w1627;
assign w1630 = ~w1628 & ~w1629;
assign w1631 = pi15 & w119;
assign w1632 = ~pi38 & pi39;
assign w1633 = ~w118 & ~w1632;
assign w1634 = pi37 & pi39;
assign w1635 = pi14 & ~w1634;
assign w1636 = ~w1633 & w1635;
assign w1637 = ~w1631 & ~w1636;
assign w1638 = pi39 & ~w1637;
assign w1639 = ~pi39 & w1637;
assign w1640 = ~w1638 & ~w1639;
assign w1641 = pi11 & w355;
assign w1642 = (pi43 & ~w353) | (pi43 & w8273) | (~w353 & w8273);
assign w1643 = pi10 & w354;
assign w1644 = ~w1641 & w8274;
assign w1645 = pi43 & w1641;
assign w1646 = ~w1644 & ~w1645;
assign w1647 = ~w1640 & ~w1646;
assign w1648 = w1640 & w1646;
assign w1649 = ~w1647 & ~w1648;
assign w1650 = pi13 & w217;
assign w1651 = (pi41 & ~w215) | (pi41 & w8275) | (~w215 & w8275);
assign w1652 = pi12 & w216;
assign w1653 = ~w1650 & w8276;
assign w1654 = pi41 & w1650;
assign w1655 = ~w1653 & ~w1654;
assign w1656 = w1649 & ~w1655;
assign w1657 = ~w1649 & w1655;
assign w1658 = ~w1656 & ~w1657;
assign w1659 = w1630 & ~w1658;
assign w1660 = ~w1630 & w1658;
assign w1661 = ~w1659 & ~w1660;
assign w1662 = w1602 & ~w1661;
assign w1663 = ~w1602 & w1661;
assign w1664 = ~w1662 & ~w1663;
assign w1665 = w1559 & ~w1664;
assign w1666 = ~w1559 & w1664;
assign w1667 = ~w1665 & ~w1666;
assign w1668 = w1558 & ~w1667;
assign w1669 = ~w1558 & w1667;
assign w1670 = ~w1668 & ~w1669;
assign w1671 = w1533 & ~w1670;
assign w1672 = ~w1533 & w1670;
assign w1673 = ~w1671 & ~w1672;
assign w1674 = ~w1528 & w1673;
assign w1675 = w1528 & ~w1673;
assign w1676 = ~w1674 & ~w1675;
assign w1677 = w1517 & ~w1676;
assign w1678 = ~w1517 & w1676;
assign w1679 = ~w1677 & ~w1678;
assign w1680 = ~w1522 & w1525;
assign w1681 = (w1679 & ~w1525) | (w1679 & w8277) | (~w1525 & w8277);
assign w1682 = w1525 & w8278;
assign w1683 = ~w1681 & ~w1682;
assign w1684 = ~w1376 & ~w1517;
assign w1685 = ~w1518 & ~w1684;
assign w1686 = w1676 & w1685;
assign w1687 = (w1557 & w1664) | (w1557 & w7555) | (w1664 & w7555);
assign w1688 = w1664 & w7556;
assign w1689 = ~w1664 & w7883;
assign w1690 = ~w1687 & ~w1688;
assign w1691 = ~w1689 & w1690;
assign w1692 = ~w1564 & ~w1596;
assign w1693 = ~pi53 & ~pi54;
assign w1694 = pi53 & pi54;
assign w1695 = ~w1693 & ~w1694;
assign w1696 = (pi55 & ~w1695) | (pi55 & w8279) | (~w1695 & w8279);
assign w1697 = w1695 & w8280;
assign w1698 = ~w1696 & ~w1697;
assign w1699 = pi02 & w1393;
assign w1700 = (pi53 & ~w1391) | (pi53 & w8281) | (~w1391 & w8281);
assign w1701 = pi01 & w1392;
assign w1702 = ~w1699 & w8282;
assign w1703 = pi53 & w1699;
assign w1704 = ~w1702 & ~w1703;
assign w1705 = w1698 & ~w1704;
assign w1706 = ~w1698 & w1704;
assign w1707 = ~w1705 & ~w1706;
assign w1708 = pi03 & ~w1260;
assign w1709 = pi04 & w1132;
assign w1710 = (pi51 & w1708) | (pi51 & w8283) | (w1708 & w8283);
assign w1711 = ~w1708 & w8284;
assign w1712 = ~w1710 & ~w1711;
assign w1713 = ~w1707 & w1712;
assign w1714 = w1707 & ~w1712;
assign w1715 = ~w1713 & ~w1714;
assign w1716 = pi55 & w1547;
assign w1717 = ~pi55 & ~w1547;
assign w1718 = ~w1716 & ~w1717;
assign w1719 = ~w1715 & w1718;
assign w1720 = w1715 & ~w1718;
assign w1721 = ~w1719 & ~w1720;
assign w1722 = w1553 & w1721;
assign w1723 = ~w1553 & ~w1721;
assign w1724 = ~w1722 & ~w1723;
assign w1725 = ~w1692 & w1724;
assign w1726 = w1692 & ~w1724;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = ~w1600 & ~w1661;
assign w1729 = ~w1601 & ~w1728;
assign w1730 = ~w1727 & ~w1729;
assign w1731 = w1727 & w1729;
assign w1732 = ~w1730 & ~w1731;
assign w1733 = (~w1591 & ~w1576) | (~w1591 & w8285) | (~w1576 & w8285);
assign w1734 = ~w1583 & ~w1733;
assign w1735 = (~w1655 & ~w1640) | (~w1655 & w8286) | (~w1640 & w8286);
assign w1736 = ~w1647 & ~w1735;
assign w1737 = w1734 & w1736;
assign w1738 = ~w1734 & ~w1736;
assign w1739 = ~w1737 & ~w1738;
assign w1740 = pi10 & w523;
assign w1741 = pi09 & ~w1570;
assign w1742 = ~w1569 & w1741;
assign w1743 = ~w1740 & ~w1742;
assign w1744 = pi45 & ~w1743;
assign w1745 = ~pi45 & w1743;
assign w1746 = ~w1744 & ~w1745;
assign w1747 = pi08 & w700;
assign w1748 = (pi47 & ~w698) | (pi47 & w8287) | (~w698 & w8287);
assign w1749 = pi07 & w699;
assign w1750 = ~w1747 & w8288;
assign w1751 = pi47 & w1747;
assign w1752 = ~w1750 & ~w1751;
assign w1753 = ~w1746 & ~w1752;
assign w1754 = w1746 & w1752;
assign w1755 = ~w1753 & ~w1754;
assign w1756 = pi06 & w909;
assign w1757 = (pi49 & ~w907) | (pi49 & w8289) | (~w907 & w8289);
assign w1758 = pi05 & w908;
assign w1759 = ~w1756 & w8290;
assign w1760 = pi49 & w1756;
assign w1761 = ~w1759 & ~w1760;
assign w1762 = w1755 & ~w1761;
assign w1763 = ~w1755 & w1761;
assign w1764 = ~w1762 & ~w1763;
assign w1765 = w1739 & ~w1764;
assign w1766 = ~w1739 & w1764;
assign w1767 = ~w1765 & ~w1766;
assign w1768 = ~w1628 & w1658;
assign w1769 = ~w1629 & ~w1768;
assign w1770 = w1767 & w1769;
assign w1771 = ~w1767 & ~w1769;
assign w1772 = ~w1770 & ~w1771;
assign w1773 = (~w1616 & ~w1618) | (~w1616 & w7557) | (~w1618 & w7557);
assign w1774 = pi18 & w56;
assign w1775 = (pi37 & ~w54) | (pi37 & w8291) | (~w54 & w8291);
assign w1776 = pi17 & w55;
assign w1777 = ~w1774 & w8292;
assign w1778 = pi37 & w1774;
assign w1779 = ~w1777 & ~w1778;
assign w1780 = pi20 & w8;
assign w1781 = (pi35 & ~w6) | (pi35 & w8293) | (~w6 & w8293);
assign w1782 = pi19 & w7;
assign w1783 = ~w1780 & w8294;
assign w1784 = pi35 & w1780;
assign w1785 = ~w1783 & ~w1784;
assign w1786 = w1779 & w1785;
assign w1787 = ~w1779 & ~w1785;
assign w1788 = ~w1786 & ~w1787;
assign w1789 = pi22 & pi32;
assign w1790 = pi21 & ~pi32;
assign w1791 = pi33 & ~w1789;
assign w1792 = ~w1790 & w1791;
assign w1793 = ~pi33 & w1789;
assign w1794 = ~w1792 & ~w1793;
assign w1795 = w1788 & ~w1794;
assign w1796 = ~w1788 & w1794;
assign w1797 = ~w1795 & ~w1796;
assign w1798 = ~w1773 & w1797;
assign w1799 = w1773 & ~w1797;
assign w1800 = ~w1798 & ~w1799;
assign w1801 = pi16 & w119;
assign w1802 = pi15 & ~w1634;
assign w1803 = ~w1633 & w1802;
assign w1804 = ~w1801 & ~w1803;
assign w1805 = pi39 & ~w1804;
assign w1806 = ~pi39 & w1804;
assign w1807 = ~w1805 & ~w1806;
assign w1808 = pi12 & w355;
assign w1809 = (pi43 & ~w353) | (pi43 & w8295) | (~w353 & w8295);
assign w1810 = pi11 & w354;
assign w1811 = ~w1808 & w8296;
assign w1812 = pi43 & w1808;
assign w1813 = ~w1811 & ~w1812;
assign w1814 = ~w1807 & ~w1813;
assign w1815 = w1807 & w1813;
assign w1816 = ~w1814 & ~w1815;
assign w1817 = pi14 & w217;
assign w1818 = (pi41 & ~w215) | (pi41 & w8297) | (~w215 & w8297);
assign w1819 = pi13 & w216;
assign w1820 = ~w1817 & w8298;
assign w1821 = pi41 & w1817;
assign w1822 = ~w1820 & ~w1821;
assign w1823 = w1816 & ~w1822;
assign w1824 = ~w1816 & w1822;
assign w1825 = ~w1823 & ~w1824;
assign w1826 = w1800 & ~w1825;
assign w1827 = ~w1800 & w1825;
assign w1828 = ~w1826 & ~w1827;
assign w1829 = w1772 & ~w1828;
assign w1830 = ~w1772 & w1828;
assign w1831 = ~w1829 & ~w1830;
assign w1832 = w1732 & ~w1831;
assign w1833 = ~w1732 & w1831;
assign w1834 = ~w1832 & ~w1833;
assign w1835 = ~w1691 & ~w1834;
assign w1836 = w1691 & w1834;
assign w1837 = ~w1835 & ~w1836;
assign w1838 = (~w1532 & w1670) | (~w1532 & w7558) | (w1670 & w7558);
assign w1839 = w1837 & ~w1838;
assign w1840 = ~w1837 & w1838;
assign w1841 = ~w1839 & ~w1840;
assign w1842 = w1686 & w1841;
assign w1843 = w1674 & w1841;
assign w1844 = ~w1674 & ~w1841;
assign w1845 = ~w1843 & ~w1844;
assign w1846 = ~w1525 & w2372;
assign w1847 = ~w1686 & ~w1845;
assign w1848 = (w1847 & w1525) | (w1847 & w8299) | (w1525 & w8299);
assign w1849 = ~w1842 & ~w1846;
assign w1850 = ~w1848 & w1849;
assign w1851 = (~w1722 & ~w1724) | (~w1722 & w8300) | (~w1724 & w8300);
assign w1852 = ~w1730 & ~w1831;
assign w1853 = ~w1852 & w7559;
assign w1854 = (~w1851 & w1852) | (~w1851 & w7560) | (w1852 & w7560);
assign w1855 = ~w1853 & ~w1854;
assign w1856 = (~w1705 & ~w1707) | (~w1705 & w7561) | (~w1707 & w7561);
assign w1857 = pi05 & w1132;
assign w1858 = pi04 & ~w1260;
assign w1859 = (pi51 & w1858) | (pi51 & w7562) | (w1858 & w7562);
assign w1860 = ~w1858 & w7563;
assign w1861 = ~w1859 & ~w1860;
assign w1862 = pi01 & w1695;
assign w1863 = ~pi54 & pi55;
assign w1864 = ~w1694 & ~w1863;
assign w1865 = pi53 & pi55;
assign w1866 = pi00 & ~w1865;
assign w1867 = ~w1864 & w1866;
assign w1868 = ~w1862 & ~w1867;
assign w1869 = pi55 & ~w1868;
assign w1870 = ~pi55 & w1868;
assign w1871 = ~w1869 & ~w1870;
assign w1872 = pi03 & w1393;
assign w1873 = (pi53 & ~w1391) | (pi53 & w8301) | (~w1391 & w8301);
assign w1874 = pi02 & w1392;
assign w1875 = ~w1872 & w8302;
assign w1876 = pi53 & w1872;
assign w1877 = ~w1875 & ~w1876;
assign w1878 = ~w1871 & ~w1877;
assign w1879 = w1871 & w1877;
assign w1880 = ~w1878 & ~w1879;
assign w1881 = w1861 & ~w1880;
assign w1882 = ~w1861 & w1880;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = w1856 & ~w1883;
assign w1885 = ~w1856 & w1883;
assign w1886 = ~w1884 & ~w1885;
assign w1887 = (~w1716 & w1715) | (~w1716 & w7564) | (w1715 & w7564);
assign w1888 = w1886 & ~w1887;
assign w1889 = ~w1886 & w1887;
assign w1890 = ~w1888 & ~w1889;
assign w1891 = ~w1737 & ~w1765;
assign w1892 = w1890 & ~w1891;
assign w1893 = ~w1890 & w1891;
assign w1894 = ~w1892 & ~w1893;
assign w1895 = ~w1770 & ~w1828;
assign w1896 = ~w1771 & ~w1895;
assign w1897 = ~w1894 & ~w1896;
assign w1898 = w1894 & w1896;
assign w1899 = ~w1897 & ~w1898;
assign w1900 = (~w1822 & ~w1807) | (~w1822 & w8303) | (~w1807 & w8303);
assign w1901 = ~w1814 & ~w1900;
assign w1902 = (~w1761 & ~w1746) | (~w1761 & w8304) | (~w1746 & w8304);
assign w1903 = ~w1753 & ~w1902;
assign w1904 = ~w1901 & ~w1903;
assign w1905 = w1901 & w1903;
assign w1906 = ~w1904 & ~w1905;
assign w1907 = pi11 & w523;
assign w1908 = pi10 & ~w1570;
assign w1909 = ~w1569 & w1908;
assign w1910 = ~w1907 & ~w1909;
assign w1911 = pi45 & ~w1910;
assign w1912 = ~pi45 & w1910;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = pi07 & w909;
assign w1915 = (pi49 & ~w907) | (pi49 & w8305) | (~w907 & w8305);
assign w1916 = pi06 & w908;
assign w1917 = ~w1914 & w8306;
assign w1918 = pi49 & w1914;
assign w1919 = ~w1917 & ~w1918;
assign w1920 = ~w1913 & ~w1919;
assign w1921 = w1913 & w1919;
assign w1922 = ~w1920 & ~w1921;
assign w1923 = pi09 & w700;
assign w1924 = (pi47 & ~w698) | (pi47 & w8307) | (~w698 & w8307);
assign w1925 = pi08 & w699;
assign w1926 = ~w1923 & w8308;
assign w1927 = pi47 & w1923;
assign w1928 = ~w1926 & ~w1927;
assign w1929 = w1922 & ~w1928;
assign w1930 = ~w1922 & w1928;
assign w1931 = ~w1929 & ~w1930;
assign w1932 = ~w1906 & ~w1931;
assign w1933 = w1906 & w1931;
assign w1934 = ~w1932 & ~w1933;
assign w1935 = ~w1798 & w1825;
assign w1936 = ~w1799 & ~w1935;
assign w1937 = w1934 & ~w1936;
assign w1938 = ~w1934 & w1936;
assign w1939 = ~w1937 & ~w1938;
assign w1940 = (~w1786 & ~w1788) | (~w1786 & w7565) | (~w1788 & w7565);
assign w1941 = pi21 & w8;
assign w1942 = (pi35 & ~w6) | (pi35 & w8309) | (~w6 & w8309);
assign w1943 = pi20 & w7;
assign w1944 = ~w1941 & w8310;
assign w1945 = pi35 & w1941;
assign w1946 = ~w1944 & ~w1945;
assign w1947 = pi19 & w56;
assign w1948 = (pi37 & ~w54) | (pi37 & w8311) | (~w54 & w8311);
assign w1949 = pi18 & w55;
assign w1950 = ~w1947 & w8312;
assign w1951 = pi37 & w1947;
assign w1952 = ~w1950 & ~w1951;
assign w1953 = w1946 & w1952;
assign w1954 = ~w1946 & ~w1952;
assign w1955 = ~w1953 & ~w1954;
assign w1956 = pi23 & pi32;
assign w1957 = pi22 & ~pi32;
assign w1958 = pi33 & ~w1956;
assign w1959 = ~w1957 & w1958;
assign w1960 = ~pi33 & w1956;
assign w1961 = ~w1959 & ~w1960;
assign w1962 = w1955 & ~w1961;
assign w1963 = ~w1955 & w1961;
assign w1964 = ~w1962 & ~w1963;
assign w1965 = ~w1940 & w1964;
assign w1966 = w1940 & ~w1964;
assign w1967 = ~w1965 & ~w1966;
assign w1968 = pi17 & w119;
assign w1969 = pi16 & ~w1634;
assign w1970 = ~w1633 & w1969;
assign w1971 = ~w1968 & ~w1970;
assign w1972 = pi39 & ~w1971;
assign w1973 = ~pi39 & w1971;
assign w1974 = ~w1972 & ~w1973;
assign w1975 = pi13 & w355;
assign w1976 = (pi43 & ~w353) | (pi43 & w8313) | (~w353 & w8313);
assign w1977 = pi12 & w354;
assign w1978 = ~w1975 & w8314;
assign w1979 = pi43 & w1975;
assign w1980 = ~w1978 & ~w1979;
assign w1981 = ~w1974 & ~w1980;
assign w1982 = w1974 & w1980;
assign w1983 = ~w1981 & ~w1982;
assign w1984 = pi15 & w217;
assign w1985 = (pi41 & ~w215) | (pi41 & w8315) | (~w215 & w8315);
assign w1986 = pi14 & w216;
assign w1987 = ~w1984 & w8316;
assign w1988 = pi41 & w1984;
assign w1989 = ~w1987 & ~w1988;
assign w1990 = w1983 & ~w1989;
assign w1991 = ~w1983 & w1989;
assign w1992 = ~w1990 & ~w1991;
assign w1993 = w1967 & w1992;
assign w1994 = ~w1967 & ~w1992;
assign w1995 = ~w1993 & ~w1994;
assign w1996 = w1939 & ~w1995;
assign w1997 = ~w1939 & w1995;
assign w1998 = ~w1996 & ~w1997;
assign w1999 = w1899 & w1998;
assign w2000 = ~w1899 & ~w1998;
assign w2001 = ~w1999 & ~w2000;
assign w2002 = ~w1855 & ~w2001;
assign w2003 = w1855 & w2001;
assign w2004 = ~w2002 & ~w2003;
assign w2005 = ~w1689 & ~w1836;
assign w2006 = w2004 & ~w2005;
assign w2007 = ~w2004 & w2005;
assign w2008 = ~w2006 & ~w2007;
assign w2009 = ~w1839 & ~w2008;
assign w2010 = w1839 & w2008;
assign w2011 = ~w2009 & ~w2010;
assign w2012 = ~w1675 & w1841;
assign w2013 = ~w1678 & w2012;
assign w2014 = ~w1842 & ~w2013;
assign w2015 = (w2014 & w1525) | (w2014 & w8317) | (w1525 & w8317);
assign w2016 = w2011 & ~w2015;
assign w2017 = ~w2011 & w2015;
assign w2018 = ~w2016 & ~w2017;
assign w2019 = (~w1854 & ~w2001) | (~w1854 & w8319) | (~w2001 & w8319);
assign w2020 = (~w1888 & ~w1890) | (~w1888 & w8320) | (~w1890 & w8320);
assign w2021 = pi57 & ~w2020;
assign w2022 = ~pi57 & w2020;
assign w2023 = ~w2021 & ~w2022;
assign w2024 = ~w1898 & ~w1998;
assign w2025 = ~w1897 & ~w2024;
assign w2026 = ~w2024 & w8321;
assign w2027 = (~w2023 & w2024) | (~w2023 & w8322) | (w2024 & w8322);
assign w2028 = ~w2026 & ~w2027;
assign w2029 = ~w1861 & ~w1879;
assign w2030 = ~pi55 & ~pi56;
assign w2031 = pi55 & pi56;
assign w2032 = ~w2030 & ~w2031;
assign w2033 = (~pi57 & ~w2032) | (~pi57 & w8323) | (~w2032 & w8323);
assign w2034 = w2032 & w8324;
assign w2035 = ~w2033 & ~w2034;
assign w2036 = (w2035 & w1871) | (w2035 & w8325) | (w1871 & w8325);
assign w2037 = ~w2029 & w2036;
assign w2038 = w1861 & ~w1878;
assign w2039 = (~w2035 & ~w1871) | (~w2035 & w8326) | (~w1871 & w8326);
assign w2040 = ~w2038 & w2039;
assign w2041 = ~w2037 & ~w2040;
assign w2042 = pi06 & w1132;
assign w2043 = pi05 & ~w1260;
assign w2044 = (pi51 & w2043) | (pi51 & w7566) | (w2043 & w7566);
assign w2045 = ~w2043 & w7567;
assign w2046 = ~w2044 & ~w2045;
assign w2047 = pi04 & w1393;
assign w2048 = ~pi52 & pi53;
assign w2049 = ~w1392 & ~w2048;
assign w2050 = pi51 & pi53;
assign w2051 = pi03 & ~w2050;
assign w2052 = ~w2049 & w2051;
assign w2053 = ~w2047 & ~w2052;
assign w2054 = pi53 & ~w2053;
assign w2055 = ~pi53 & w2053;
assign w2056 = ~w2054 & ~w2055;
assign w2057 = pi02 & w1695;
assign w2058 = (pi55 & ~w1693) | (pi55 & w8327) | (~w1693 & w8327);
assign w2059 = pi01 & w1694;
assign w2060 = ~w2057 & w8328;
assign w2061 = pi55 & w2057;
assign w2062 = ~w2060 & ~w2061;
assign w2063 = ~w2056 & ~w2062;
assign w2064 = w2056 & w2062;
assign w2065 = ~w2063 & ~w2064;
assign w2066 = w2046 & ~w2065;
assign w2067 = ~w2046 & w2065;
assign w2068 = ~w2066 & ~w2067;
assign w2069 = w2041 & w2068;
assign w2070 = ~w2041 & ~w2068;
assign w2071 = ~w2069 & ~w2070;
assign w2072 = ~w1884 & w2071;
assign w2073 = w1884 & ~w2071;
assign w2074 = ~w2072 & ~w2073;
assign w2075 = ~w1904 & ~w1933;
assign w2076 = w2074 & ~w2075;
assign w2077 = ~w2074 & w2075;
assign w2078 = ~w2076 & ~w2077;
assign w2079 = ~w1938 & w1995;
assign w2080 = ~w1937 & ~w2079;
assign w2081 = w2078 & ~w2080;
assign w2082 = ~w2078 & w2080;
assign w2083 = ~w2081 & ~w2082;
assign w2084 = (~w1989 & ~w1974) | (~w1989 & w8329) | (~w1974 & w8329);
assign w2085 = ~w1981 & ~w2084;
assign w2086 = (~w1928 & ~w1913) | (~w1928 & w8330) | (~w1913 & w8330);
assign w2087 = ~w1920 & ~w2086;
assign w2088 = w2085 & w2087;
assign w2089 = ~w2085 & ~w2087;
assign w2090 = ~w2088 & ~w2089;
assign w2091 = pi11 & ~w612;
assign w2092 = pi12 & w523;
assign w2093 = (pi45 & w2091) | (pi45 & w7568) | (w2091 & w7568);
assign w2094 = ~w2091 & w7569;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = pi10 & w700;
assign w2097 = ~pi46 & pi47;
assign w2098 = ~w699 & ~w2097;
assign w2099 = pi45 & pi47;
assign w2100 = pi09 & ~w2099;
assign w2101 = ~w2098 & w2100;
assign w2102 = ~w2096 & ~w2101;
assign w2103 = pi47 & ~w2102;
assign w2104 = ~pi47 & w2102;
assign w2105 = ~w2103 & ~w2104;
assign w2106 = pi08 & w909;
assign w2107 = (pi49 & ~w907) | (pi49 & w8331) | (~w907 & w8331);
assign w2108 = pi07 & w908;
assign w2109 = ~w2106 & w8332;
assign w2110 = pi49 & w2106;
assign w2111 = ~w2109 & ~w2110;
assign w2112 = ~w2105 & ~w2111;
assign w2113 = w2105 & w2111;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = w2095 & ~w2114;
assign w2116 = ~w2095 & w2114;
assign w2117 = ~w2115 & ~w2116;
assign w2118 = ~w2090 & w2117;
assign w2119 = w2090 & ~w2117;
assign w2120 = ~w2118 & ~w2119;
assign w2121 = ~w1966 & ~w1992;
assign w2122 = ~w1965 & ~w2121;
assign w2123 = w2120 & ~w2122;
assign w2124 = ~w2120 & w2122;
assign w2125 = ~w2123 & ~w2124;
assign w2126 = (~w1953 & ~w1955) | (~w1953 & w7570) | (~w1955 & w7570);
assign w2127 = pi17 & ~w167;
assign w2128 = pi18 & w119;
assign w2129 = (pi39 & w2127) | (pi39 & w7571) | (w2127 & w7571);
assign w2130 = ~w2127 & w7572;
assign w2131 = ~w2129 & ~w2130;
assign w2132 = pi16 & w217;
assign w2133 = pi15 & ~w802;
assign w2134 = ~w801 & w2133;
assign w2135 = ~w2132 & ~w2134;
assign w2136 = pi41 & ~w2135;
assign w2137 = ~pi41 & w2135;
assign w2138 = ~w2136 & ~w2137;
assign w2139 = pi14 & w355;
assign w2140 = (pi43 & ~w353) | (pi43 & w8333) | (~w353 & w8333);
assign w2141 = pi13 & w354;
assign w2142 = ~w2139 & w8334;
assign w2143 = pi43 & w2139;
assign w2144 = ~w2142 & ~w2143;
assign w2145 = ~w2138 & ~w2144;
assign w2146 = w2138 & w2144;
assign w2147 = ~w2145 & ~w2146;
assign w2148 = w2131 & ~w2147;
assign w2149 = ~w2131 & w2147;
assign w2150 = ~w2148 & ~w2149;
assign w2151 = w2126 & w2150;
assign w2152 = ~w2126 & ~w2150;
assign w2153 = ~w2151 & ~w2152;
assign w2154 = pi21 & ~w25;
assign w2155 = pi22 & w8;
assign w2156 = (pi35 & w2154) | (pi35 & w8335) | (w2154 & w8335);
assign w2157 = ~w2154 & w8336;
assign w2158 = ~w2156 & ~w2157;
assign w2159 = pi20 & w56;
assign w2160 = (pi37 & ~w54) | (pi37 & w8337) | (~w54 & w8337);
assign w2161 = pi19 & w55;
assign w2162 = ~w2159 & w8338;
assign w2163 = pi37 & w2159;
assign w2164 = pi24 & pi32;
assign w2165 = pi23 & ~pi32;
assign w2166 = pi33 & ~w2164;
assign w2167 = ~w2165 & w2166;
assign w2168 = ~pi33 & w2164;
assign w2169 = ~w2167 & ~w2168;
assign w2170 = (w2169 & w2162) | (w2169 & w7573) | (w2162 & w7573);
assign w2171 = ~w2162 & w7574;
assign w2172 = ~w2170 & ~w2171;
assign w2173 = w2158 & w2172;
assign w2174 = ~w2158 & ~w2172;
assign w2175 = ~w2173 & ~w2174;
assign w2176 = w2153 & ~w2175;
assign w2177 = ~w2153 & w2175;
assign w2178 = ~w2176 & ~w2177;
assign w2179 = w2125 & ~w2178;
assign w2180 = ~w2125 & w2178;
assign w2181 = ~w2179 & ~w2180;
assign w2182 = w2083 & w2181;
assign w2183 = ~w2083 & ~w2181;
assign w2184 = ~w2182 & ~w2183;
assign w2185 = w2028 & ~w2184;
assign w2186 = ~w2028 & w2184;
assign w2187 = ~w2185 & ~w2186;
assign w2188 = w2019 & w2187;
assign w2189 = ~w2019 & ~w2187;
assign w2190 = ~w2188 & ~w2189;
assign w2191 = ~w2006 & w2190;
assign w2192 = w2006 & ~w2190;
assign w2193 = ~w2191 & ~w2192;
assign w2194 = (w2015 & w8339) | (w2015 & w8340) | (w8339 & w8340);
assign w2195 = ~w2193 & w9079;
assign w2196 = ~w2194 & ~w2195;
assign w2197 = (~w2072 & ~w2074) | (~w2072 & w8341) | (~w2074 & w8341);
assign w2198 = ~w2082 & ~w2181;
assign w2199 = (~w2197 & w2198) | (~w2197 & w7575) | (w2198 & w7575);
assign w2200 = ~w2198 & w7576;
assign w2201 = ~w2199 & ~w2200;
assign w2202 = ~w2046 & ~w2064;
assign w2203 = pi01 & w2032;
assign w2204 = pi57 & w2030;
assign w2205 = ~pi57 & w2031;
assign w2206 = ~w2204 & ~w2205;
assign w2207 = pi00 & ~w2206;
assign w2208 = (pi57 & w2207) | (pi57 & w7577) | (w2207 & w7577);
assign w2209 = ~w2207 & w7578;
assign w2210 = ~w2208 & ~w2209;
assign w2211 = ~w2063 & w2210;
assign w2212 = ~w2202 & w2211;
assign w2213 = w2046 & ~w2063;
assign w2214 = ~w2064 & ~w2210;
assign w2215 = ~w2213 & w2214;
assign w2216 = ~w2212 & ~w2215;
assign w2217 = pi06 & ~w1260;
assign w2218 = pi07 & w1132;
assign w2219 = (pi51 & w2217) | (pi51 & w7579) | (w2217 & w7579);
assign w2220 = ~w2217 & w7580;
assign w2221 = ~w2219 & ~w2220;
assign w2222 = pi05 & w1393;
assign w2223 = pi04 & ~w2050;
assign w2224 = ~w2049 & w2223;
assign w2225 = ~w2222 & ~w2224;
assign w2226 = pi53 & ~w2225;
assign w2227 = ~pi53 & w2225;
assign w2228 = ~w2226 & ~w2227;
assign w2229 = pi03 & w1695;
assign w2230 = (pi55 & ~w1693) | (pi55 & w8342) | (~w1693 & w8342);
assign w2231 = pi02 & w1694;
assign w2232 = ~w2229 & w8343;
assign w2233 = pi55 & w2229;
assign w2234 = ~w2232 & ~w2233;
assign w2235 = ~w2228 & ~w2234;
assign w2236 = w2228 & w2234;
assign w2237 = ~w2235 & ~w2236;
assign w2238 = w2221 & ~w2237;
assign w2239 = ~w2221 & w2237;
assign w2240 = ~w2238 & ~w2239;
assign w2241 = ~w2216 & w2240;
assign w2242 = w2216 & ~w2240;
assign w2243 = ~w2241 & ~w2242;
assign w2244 = ~w2040 & ~w2069;
assign w2245 = w2243 & w2244;
assign w2246 = ~w2243 & ~w2244;
assign w2247 = ~w2245 & ~w2246;
assign w2248 = ~w2088 & ~w2119;
assign w2249 = ~w2247 & w2248;
assign w2250 = w2247 & ~w2248;
assign w2251 = ~w2249 & ~w2250;
assign w2252 = (~w2124 & ~w2178) | (~w2124 & w8344) | (~w2178 & w8344);
assign w2253 = ~w2251 & ~w2252;
assign w2254 = w2251 & w2252;
assign w2255 = ~w2253 & ~w2254;
assign w2256 = (w2175 & ~w2150) | (w2175 & w7581) | (~w2150 & w7581);
assign w2257 = ~w2152 & ~w2256;
assign w2258 = ~w2131 & ~w2146;
assign w2259 = ~w2145 & ~w2258;
assign w2260 = ~w2095 & ~w2113;
assign w2261 = ~w2112 & ~w2260;
assign w2262 = ~w2259 & ~w2261;
assign w2263 = w2259 & w2261;
assign w2264 = ~w2262 & ~w2263;
assign w2265 = pi12 & ~w612;
assign w2266 = pi13 & w523;
assign w2267 = (pi45 & w2265) | (pi45 & w7582) | (w2265 & w7582);
assign w2268 = ~w2265 & w7583;
assign w2269 = ~w2267 & ~w2268;
assign w2270 = pi09 & w909;
assign w2271 = ~pi48 & pi49;
assign w2272 = ~w908 & ~w2271;
assign w2273 = pi47 & pi49;
assign w2274 = pi08 & ~w2273;
assign w2275 = ~w2272 & w2274;
assign w2276 = ~w2270 & ~w2275;
assign w2277 = pi49 & ~w2276;
assign w2278 = ~pi49 & w2276;
assign w2279 = ~w2277 & ~w2278;
assign w2280 = pi11 & w700;
assign w2281 = pi10 & ~w2099;
assign w2282 = ~w2098 & w2281;
assign w2283 = ~w2280 & ~w2282;
assign w2284 = pi47 & ~w2283;
assign w2285 = ~pi47 & w2283;
assign w2286 = ~w2284 & ~w2285;
assign w2287 = ~w2279 & ~w2286;
assign w2288 = w2279 & w2286;
assign w2289 = ~w2287 & ~w2288;
assign w2290 = w2269 & ~w2289;
assign w2291 = ~w2269 & w2289;
assign w2292 = ~w2290 & ~w2291;
assign w2293 = w2264 & ~w2292;
assign w2294 = ~w2264 & w2292;
assign w2295 = ~w2293 & ~w2294;
assign w2296 = w2257 & ~w2295;
assign w2297 = ~w2257 & w2295;
assign w2298 = ~w2296 & ~w2297;
assign w2299 = (~w2171 & ~w2172) | (~w2171 & w8345) | (~w2172 & w8345);
assign w2300 = pi18 & ~w167;
assign w2301 = pi19 & w119;
assign w2302 = (pi39 & w2300) | (pi39 & w7584) | (w2300 & w7584);
assign w2303 = ~w2300 & w7585;
assign w2304 = ~w2302 & ~w2303;
assign w2305 = pi17 & w217;
assign w2306 = pi16 & ~w802;
assign w2307 = ~w801 & w2306;
assign w2308 = ~w2305 & ~w2307;
assign w2309 = pi41 & ~w2308;
assign w2310 = ~pi41 & w2308;
assign w2311 = ~w2309 & ~w2310;
assign w2312 = pi15 & w355;
assign w2313 = (pi43 & ~w353) | (pi43 & w8346) | (~w353 & w8346);
assign w2314 = pi14 & w354;
assign w2315 = ~w2312 & w8347;
assign w2316 = pi43 & w2312;
assign w2317 = ~w2315 & ~w2316;
assign w2318 = ~w2311 & ~w2317;
assign w2319 = w2311 & w2317;
assign w2320 = ~w2318 & ~w2319;
assign w2321 = w2304 & ~w2320;
assign w2322 = ~w2304 & w2320;
assign w2323 = ~w2321 & ~w2322;
assign w2324 = w2299 & w2323;
assign w2325 = ~w2299 & ~w2323;
assign w2326 = ~w2324 & ~w2325;
assign w2327 = pi22 & ~w25;
assign w2328 = (pi35 & w2327) | (pi35 & w7586) | (w2327 & w7586);
assign w2329 = ~w2327 & w7587;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = pi37 & w54;
assign w2332 = ~w90 & ~w2331;
assign w2333 = pi20 & ~w2332;
assign w2334 = (pi37 & w2333) | (pi37 & w7588) | (w2333 & w7588);
assign w2335 = ~w2333 & w7589;
assign w2336 = ~w2334 & ~w2335;
assign w2337 = w2330 & w2336;
assign w2338 = ~w2330 & ~w2336;
assign w2339 = ~w2337 & ~w2338;
assign w2340 = pi25 & pi32;
assign w2341 = pi24 & ~pi32;
assign w2342 = pi33 & ~w2340;
assign w2343 = ~w2341 & w2342;
assign w2344 = ~pi33 & w2340;
assign w2345 = ~w2343 & ~w2344;
assign w2346 = w2339 & ~w2345;
assign w2347 = ~w2339 & w2345;
assign w2348 = ~w2346 & ~w2347;
assign w2349 = w2326 & w2348;
assign w2350 = ~w2326 & ~w2348;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = w2298 & ~w2351;
assign w2353 = ~w2298 & w2351;
assign w2354 = ~w2352 & ~w2353;
assign w2355 = w2255 & ~w2354;
assign w2356 = ~w2255 & w2354;
assign w2357 = ~w2355 & ~w2356;
assign w2358 = ~w2201 & ~w2357;
assign w2359 = w2201 & w2357;
assign w2360 = ~w2358 & ~w2359;
assign w2361 = ~w2027 & w2184;
assign w2362 = (~w2021 & ~w2025) | (~w2021 & w7590) | (~w2025 & w7590);
assign w2363 = ~w2361 & w2362;
assign w2364 = w2184 & w8348;
assign w2365 = ~w2363 & ~w2364;
assign w2366 = w2360 & ~w2365;
assign w2367 = ~w2360 & w2365;
assign w2368 = ~w2366 & ~w2367;
assign w2369 = w2189 & ~w2368;
assign w2370 = ~w2189 & w2368;
assign w2371 = ~w2369 & ~w2370;
assign w2372 = ~w1679 & w1845;
assign w2373 = ~w1679 & w7884;
assign w2374 = ~w1247 & w2373;
assign w2375 = w1524 & w2372;
assign w2376 = (~w2006 & ~w2008) | (~w2006 & w7885) | (~w2008 & w7885);
assign w2377 = w2190 & ~w2376;
assign w2378 = w2014 & ~w2377;
assign w2379 = ~w2375 & w2378;
assign w2380 = ~w2374 & w2379;
assign w2381 = w2011 & ~w2193;
assign w2382 = (~w2377 & w2193) | (~w2377 & w7886) | (w2193 & w7886);
assign w2383 = (~w2382 & ~w2379) | (~w2382 & w7887) | (~w2379 & w7887);
assign w2384 = w2371 & w2383;
assign w2385 = ~w2371 & ~w2383;
assign w2386 = ~w2384 & ~w2385;
assign w2387 = ~w2200 & ~w2359;
assign w2388 = ~pi57 & ~pi58;
assign w2389 = pi57 & pi58;
assign w2390 = ~w2388 & ~w2389;
assign w2391 = pi00 & w2390;
assign w2392 = (~w2245 & ~w2247) | (~w2245 & w8349) | (~w2247 & w8349);
assign w2393 = w2391 & ~w2392;
assign w2394 = ~w2391 & w2392;
assign w2395 = ~w2393 & ~w2394;
assign w2396 = ~w2254 & w2354;
assign w2397 = ~w2253 & ~w2396;
assign w2398 = (~w2395 & w2396) | (~w2395 & w8350) | (w2396 & w8350);
assign w2399 = ~w2396 & w8351;
assign w2400 = ~w2398 & ~w2399;
assign w2401 = ~w2212 & ~w2242;
assign w2402 = ~w2263 & w2292;
assign w2403 = ~w2262 & ~w2402;
assign w2404 = w2401 & ~w2403;
assign w2405 = ~w2401 & w2403;
assign w2406 = ~w2404 & ~w2405;
assign w2407 = pi01 & ~w2206;
assign w2408 = pi02 & w2032;
assign w2409 = (pi57 & w2407) | (pi57 & w8352) | (w2407 & w8352);
assign w2410 = ~w2407 & w8353;
assign w2411 = ~w2409 & ~w2410;
assign w2412 = ~w2221 & ~w2236;
assign w2413 = ~w2412 & w7591;
assign w2414 = (~w2411 & w2412) | (~w2411 & w8354) | (w2412 & w8354);
assign w2415 = ~w2413 & ~w2414;
assign w2416 = pi08 & w1132;
assign w2417 = ~pi50 & pi51;
assign w2418 = ~w1131 & ~w2417;
assign w2419 = pi49 & pi51;
assign w2420 = pi07 & ~w2419;
assign w2421 = ~w2418 & w2420;
assign w2422 = ~w2416 & ~w2421;
assign w2423 = pi51 & ~w2422;
assign w2424 = ~pi51 & w2422;
assign w2425 = ~w2423 & ~w2424;
assign w2426 = pi04 & w1695;
assign w2427 = (pi55 & ~w1693) | (pi55 & w7592) | (~w1693 & w7592);
assign w2428 = ~pi55 & w1694;
assign w2429 = w1694 & w8355;
assign w2430 = ~w2426 & w8356;
assign w2431 = w1695 & w9010;
assign w2432 = ~w2430 & ~w2431;
assign w2433 = ~w2425 & ~w2432;
assign w2434 = w2425 & w2432;
assign w2435 = ~w2433 & ~w2434;
assign w2436 = pi06 & w1393;
assign w2437 = (pi53 & ~w1391) | (pi53 & w8357) | (~w1391 & w8357);
assign w2438 = w1392 & w9011;
assign w2439 = ~w2436 & ~w2437;
assign w2440 = w1393 & w8358;
assign w2441 = (~w2440 & ~w2439) | (~w2440 & w8359) | (~w2439 & w8359);
assign w2442 = w2435 & ~w2441;
assign w2443 = ~w2435 & w2441;
assign w2444 = ~w2442 & ~w2443;
assign w2445 = w2415 & ~w2444;
assign w2446 = ~w2415 & w2444;
assign w2447 = ~w2445 & ~w2446;
assign w2448 = w2406 & ~w2447;
assign w2449 = ~w2406 & w2447;
assign w2450 = ~w2448 & ~w2449;
assign w2451 = ~w2297 & ~w2351;
assign w2452 = ~w2296 & ~w2451;
assign w2453 = w2450 & ~w2452;
assign w2454 = ~w2450 & w2452;
assign w2455 = ~w2453 & ~w2454;
assign w2456 = ~w2269 & ~w2288;
assign w2457 = ~w2287 & ~w2456;
assign w2458 = ~w2304 & ~w2319;
assign w2459 = ~w2318 & ~w2458;
assign w2460 = w2457 & w2459;
assign w2461 = ~w2457 & ~w2459;
assign w2462 = ~w2460 & ~w2461;
assign w2463 = pi14 & w523;
assign w2464 = pi13 & ~w1570;
assign w2465 = ~w1569 & w2464;
assign w2466 = ~w2463 & ~w2465;
assign w2467 = pi45 & ~w2466;
assign w2468 = ~pi45 & w2466;
assign w2469 = ~w2467 & ~w2468;
assign w2470 = pi12 & w700;
assign w2471 = (pi47 & ~w698) | (pi47 & w7593) | (~w698 & w7593);
assign w2472 = w699 & w8360;
assign w2473 = ~w2470 & w8361;
assign w2474 = w700 & w9012;
assign w2475 = ~w2473 & ~w2474;
assign w2476 = ~w2469 & ~w2475;
assign w2477 = w2469 & w2475;
assign w2478 = ~w2476 & ~w2477;
assign w2479 = pi10 & w909;
assign w2480 = (pi49 & ~w907) | (pi49 & w8362) | (~w907 & w8362);
assign w2481 = ~pi49 & w908;
assign w2482 = w908 & w8363;
assign w2483 = ~w2479 & w8364;
assign w2484 = w909 & w9013;
assign w2485 = ~w2483 & ~w2484;
assign w2486 = w2478 & ~w2485;
assign w2487 = ~w2478 & w2485;
assign w2488 = ~w2486 & ~w2487;
assign w2489 = w2462 & ~w2488;
assign w2490 = ~w2462 & w2488;
assign w2491 = ~w2489 & ~w2490;
assign w2492 = ~w2325 & ~w2348;
assign w2493 = ~w2324 & ~w2492;
assign w2494 = ~w2491 & ~w2493;
assign w2495 = w2491 & w2493;
assign w2496 = ~w2494 & ~w2495;
assign w2497 = ~w2338 & ~w2345;
assign w2498 = ~w2337 & ~w2497;
assign w2499 = pi20 & w119;
assign w2500 = pi19 & ~w1634;
assign w2501 = ~w1633 & w2500;
assign w2502 = ~w2499 & ~w2501;
assign w2503 = pi39 & ~w2502;
assign w2504 = ~pi39 & w2502;
assign w2505 = ~w2503 & ~w2504;
assign w2506 = pi18 & w217;
assign w2507 = (pi41 & ~w215) | (pi41 & w7594) | (~w215 & w7594);
assign w2508 = w216 & w8365;
assign w2509 = ~w2506 & w8366;
assign w2510 = w217 & w9014;
assign w2511 = ~w2509 & ~w2510;
assign w2512 = ~w2505 & ~w2511;
assign w2513 = w2505 & w2511;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = pi16 & w355;
assign w2516 = (pi43 & ~w353) | (pi43 & w8367) | (~w353 & w8367);
assign w2517 = w438 & w9015;
assign w2518 = ~w2515 & ~w2516;
assign w2519 = w355 & w8368;
assign w2520 = (~w2519 & ~w2518) | (~w2519 & w8369) | (~w2518 & w8369);
assign w2521 = w2514 & ~w2520;
assign w2522 = ~w2514 & w2520;
assign w2523 = ~w2521 & ~w2522;
assign w2524 = ~w2498 & ~w2523;
assign w2525 = w2498 & w2523;
assign w2526 = ~w2524 & ~w2525;
assign w2527 = pi22 & w56;
assign w2528 = (pi37 & ~w54) | (pi37 & w7595) | (~w54 & w7595);
assign w2529 = w55 & w8370;
assign w2530 = ~w2527 & w8371;
assign w2531 = w56 & w9016;
assign w2532 = ~w2530 & ~w2531;
assign w2533 = pi24 & w8;
assign w2534 = (pi35 & ~w6) | (pi35 & w7596) | (~w6 & w7596);
assign w2535 = w7 & w8372;
assign w2536 = ~w2533 & w8373;
assign w2537 = w8 & w9017;
assign w2538 = ~w2536 & ~w2537;
assign w2539 = w2532 & w2538;
assign w2540 = ~w2532 & ~w2538;
assign w2541 = ~w2539 & ~w2540;
assign w2542 = pi26 & pi32;
assign w2543 = pi25 & ~pi32;
assign w2544 = pi33 & ~w2542;
assign w2545 = ~w2543 & w2544;
assign w2546 = ~pi33 & w2542;
assign w2547 = ~w2545 & ~w2546;
assign w2548 = w2541 & ~w2547;
assign w2549 = ~w2541 & w2547;
assign w2550 = ~w2548 & ~w2549;
assign w2551 = w2526 & ~w2550;
assign w2552 = ~w2526 & w2550;
assign w2553 = ~w2551 & ~w2552;
assign w2554 = w2496 & ~w2553;
assign w2555 = ~w2496 & w2553;
assign w2556 = ~w2554 & ~w2555;
assign w2557 = w2455 & w2556;
assign w2558 = ~w2455 & ~w2556;
assign w2559 = ~w2557 & ~w2558;
assign w2560 = ~w2400 & ~w2559;
assign w2561 = w2400 & w2559;
assign w2562 = ~w2560 & ~w2561;
assign w2563 = ~w2387 & w2562;
assign w2564 = w2387 & ~w2562;
assign w2565 = ~w2563 & ~w2564;
assign w2566 = (~w2363 & ~w2365) | (~w2363 & w7597) | (~w2365 & w7597);
assign w2567 = ~w2565 & ~w2566;
assign w2568 = w2565 & w2566;
assign w2569 = ~w2567 & ~w2568;
assign w2570 = ~w2189 & w2376;
assign w2571 = ~w2188 & ~w2368;
assign w2572 = ~w2570 & w2571;
assign w2573 = (w2383 & w8374) | (w2383 & w8375) | (w8374 & w8375);
assign w2574 = ~w2569 & w9080;
assign w2575 = ~w2573 & ~w2574;
assign w2576 = ~w2568 & ~w2573;
assign w2577 = w2393 & ~w2559;
assign w2578 = (w2393 & w2396) | (w2393 & w7598) | (w2396 & w7598);
assign w2579 = (~w2393 & w2397) | (~w2393 & w7599) | (w2397 & w7599);
assign w2580 = w2559 & w2579;
assign w2581 = ~w2399 & ~w2578;
assign w2582 = ~w2577 & w2581;
assign w2583 = ~w2580 & w2582;
assign w2584 = (~w2404 & ~w2406) | (~w2404 & w8376) | (~w2406 & w8376);
assign w2585 = w2390 & w8377;
assign w2586 = pi59 & w2388;
assign w2587 = ~pi59 & w2389;
assign w2588 = ~w2586 & ~w2587;
assign w2589 = pi00 & ~w2588;
assign w2590 = pi01 & w2390;
assign w2591 = (w2585 & w2589) | (w2585 & w8378) | (w2589 & w8378);
assign w2592 = ~w2589 & w8379;
assign w2593 = ~w2591 & ~w2592;
assign w2594 = w2584 & w2593;
assign w2595 = ~w2584 & ~w2593;
assign w2596 = ~w2594 & ~w2595;
assign w2597 = ~w2454 & ~w2556;
assign w2598 = ~w2453 & ~w2597;
assign w2599 = ~w2597 & w8380;
assign w2600 = (~w2596 & w2597) | (~w2596 & w8381) | (w2597 & w8381);
assign w2601 = ~w2599 & ~w2600;
assign w2602 = (~w2414 & ~w2444) | (~w2414 & w8382) | (~w2444 & w8382);
assign w2603 = ~w2460 & w2488;
assign w2604 = ~w2461 & ~w2603;
assign w2605 = w2602 & w2604;
assign w2606 = ~w2602 & ~w2604;
assign w2607 = ~w2605 & ~w2606;
assign w2608 = pi02 & ~w2206;
assign w2609 = pi03 & w2032;
assign w2610 = (pi57 & w2608) | (pi57 & w8383) | (w2608 & w8383);
assign w2611 = ~w2608 & w8384;
assign w2612 = ~w2610 & ~w2611;
assign w2613 = (~w2441 & ~w2425) | (~w2441 & w8385) | (~w2425 & w8385);
assign w2614 = ~w2433 & ~w2613;
assign w2615 = ~w2613 & w7600;
assign w2616 = ~w2612 & ~w2614;
assign w2617 = ~w2615 & ~w2616;
assign w2618 = pi09 & w1132;
assign w2619 = pi08 & ~w2419;
assign w2620 = ~w2418 & w2619;
assign w2621 = ~w2618 & ~w2620;
assign w2622 = pi51 & ~w2621;
assign w2623 = ~pi51 & w2621;
assign w2624 = ~w2622 & ~w2623;
assign w2625 = pi05 & w1695;
assign w2626 = (pi55 & ~w1693) | (pi55 & w7601) | (~w1693 & w7601);
assign w2627 = w1694 & w8386;
assign w2628 = ~w2625 & w8387;
assign w2629 = w1695 & w9018;
assign w2630 = ~w2628 & ~w2629;
assign w2631 = ~w2624 & ~w2630;
assign w2632 = w2624 & w2630;
assign w2633 = ~w2631 & ~w2632;
assign w2634 = pi07 & w1393;
assign w2635 = (pi53 & ~w1391) | (pi53 & w8388) | (~w1391 & w8388);
assign w2636 = w1392 & w9019;
assign w2637 = ~w2634 & ~w2635;
assign w2638 = w1393 & w8389;
assign w2639 = (~w2638 & ~w2637) | (~w2638 & w8390) | (~w2637 & w8390);
assign w2640 = w2633 & ~w2639;
assign w2641 = ~w2633 & w2639;
assign w2642 = ~w2640 & ~w2641;
assign w2643 = w2617 & ~w2642;
assign w2644 = ~w2617 & w2642;
assign w2645 = ~w2643 & ~w2644;
assign w2646 = ~w2607 & ~w2645;
assign w2647 = w2607 & w2645;
assign w2648 = ~w2646 & ~w2647;
assign w2649 = ~w2495 & w2553;
assign w2650 = ~w2494 & ~w2649;
assign w2651 = w2648 & w2650;
assign w2652 = ~w2648 & ~w2650;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = (w2550 & ~w2523) | (w2550 & w8391) | (~w2523 & w8391);
assign w2655 = ~w2524 & ~w2654;
assign w2656 = (~w2520 & ~w2505) | (~w2520 & w8392) | (~w2505 & w8392);
assign w2657 = ~w2512 & ~w2656;
assign w2658 = (~w2485 & ~w2469) | (~w2485 & w8393) | (~w2469 & w8393);
assign w2659 = ~w2476 & ~w2658;
assign w2660 = ~w2657 & ~w2659;
assign w2661 = w2657 & w2659;
assign w2662 = ~w2660 & ~w2661;
assign w2663 = pi15 & w523;
assign w2664 = pi14 & ~w1570;
assign w2665 = ~w1569 & w2664;
assign w2666 = ~w2663 & ~w2665;
assign w2667 = pi45 & ~w2666;
assign w2668 = ~pi45 & w2666;
assign w2669 = ~w2667 & ~w2668;
assign w2670 = pi11 & w909;
assign w2671 = (pi49 & ~w907) | (pi49 & w7602) | (~w907 & w7602);
assign w2672 = w908 & w8394;
assign w2673 = ~w2670 & w8395;
assign w2674 = w909 & w9020;
assign w2675 = ~w2673 & ~w2674;
assign w2676 = ~w2669 & ~w2675;
assign w2677 = w2669 & w2675;
assign w2678 = ~w2676 & ~w2677;
assign w2679 = pi13 & w700;
assign w2680 = (pi47 & ~w698) | (pi47 & w8396) | (~w698 & w8396);
assign w2681 = w699 & w9021;
assign w2682 = ~w2679 & ~w2680;
assign w2683 = w700 & w8397;
assign w2684 = (~w2683 & ~w2682) | (~w2683 & w8398) | (~w2682 & w8398);
assign w2685 = w2678 & ~w2684;
assign w2686 = ~w2678 & w2684;
assign w2687 = ~w2685 & ~w2686;
assign w2688 = w2662 & ~w2687;
assign w2689 = ~w2662 & w2687;
assign w2690 = ~w2688 & ~w2689;
assign w2691 = w2655 & ~w2690;
assign w2692 = ~w2655 & w2690;
assign w2693 = ~w2691 & ~w2692;
assign w2694 = (~w2539 & ~w2541) | (~w2539 & w7603) | (~w2541 & w7603);
assign w2695 = pi23 & w56;
assign w2696 = (pi37 & ~w54) | (pi37 & w8399) | (~w54 & w8399);
assign w2697 = pi22 & w55;
assign w2698 = ~w2695 & w8400;
assign w2699 = w56 & w9022;
assign w2700 = ~w2698 & ~w2699;
assign w2701 = pi25 & w8;
assign w2702 = (pi35 & ~w6) | (pi35 & w8401) | (~w6 & w8401);
assign w2703 = pi24 & w7;
assign w2704 = ~w2701 & w8402;
assign w2705 = w8 & w9023;
assign w2706 = ~w2704 & ~w2705;
assign w2707 = w2700 & w2706;
assign w2708 = ~w2700 & ~w2706;
assign w2709 = ~w2707 & ~w2708;
assign w2710 = pi27 & pi32;
assign w2711 = pi26 & ~pi32;
assign w2712 = pi33 & ~w2710;
assign w2713 = ~w2711 & w2712;
assign w2714 = ~pi33 & w2710;
assign w2715 = ~w2713 & ~w2714;
assign w2716 = w2709 & ~w2715;
assign w2717 = ~w2709 & w2715;
assign w2718 = ~w2716 & ~w2717;
assign w2719 = ~w2694 & w2718;
assign w2720 = w2694 & ~w2718;
assign w2721 = ~w2719 & ~w2720;
assign w2722 = pi21 & w119;
assign w2723 = pi20 & ~w1634;
assign w2724 = ~w1633 & w2723;
assign w2725 = ~w2722 & ~w2724;
assign w2726 = pi39 & ~w2725;
assign w2727 = ~pi39 & w2725;
assign w2728 = ~w2726 & ~w2727;
assign w2729 = pi17 & w355;
assign w2730 = (pi43 & ~w353) | (pi43 & w7604) | (~w353 & w7604);
assign w2731 = w438 & w8403;
assign w2732 = ~w2729 & w8404;
assign w2733 = w355 & w9024;
assign w2734 = ~w2732 & ~w2733;
assign w2735 = ~w2728 & ~w2734;
assign w2736 = w2728 & w2734;
assign w2737 = ~w2735 & ~w2736;
assign w2738 = pi19 & w217;
assign w2739 = (pi41 & ~w215) | (pi41 & w8405) | (~w215 & w8405);
assign w2740 = w216 & w9025;
assign w2741 = ~w2738 & ~w2739;
assign w2742 = w217 & w8406;
assign w2743 = (~w2742 & ~w2741) | (~w2742 & w8407) | (~w2741 & w8407);
assign w2744 = w2737 & ~w2743;
assign w2745 = ~w2737 & w2743;
assign w2746 = ~w2744 & ~w2745;
assign w2747 = w2721 & ~w2746;
assign w2748 = ~w2721 & w2746;
assign w2749 = ~w2747 & ~w2748;
assign w2750 = w2693 & ~w2749;
assign w2751 = ~w2693 & w2749;
assign w2752 = ~w2750 & ~w2751;
assign w2753 = w2653 & ~w2752;
assign w2754 = ~w2653 & w2752;
assign w2755 = ~w2753 & ~w2754;
assign w2756 = w2601 & w2755;
assign w2757 = ~w2601 & ~w2755;
assign w2758 = ~w2756 & ~w2757;
assign w2759 = ~w2583 & w2758;
assign w2760 = w2583 & ~w2758;
assign w2761 = ~w2759 & ~w2760;
assign w2762 = w2563 & w2761;
assign w2763 = ~w2563 & ~w2761;
assign w2764 = ~w2762 & ~w2763;
assign w2765 = w2576 & w2764;
assign w2766 = ~w2576 & ~w2764;
assign w2767 = ~w2765 & ~w2766;
assign w2768 = w2393 & w2561;
assign w2769 = (~w2768 & w2583) | (~w2768 & w8408) | (w2583 & w8408);
assign w2770 = (w2595 & w2597) | (w2595 & w8409) | (w2597 & w8409);
assign w2771 = ~w2597 & w7605;
assign w2772 = w2755 & w2771;
assign w2773 = (~w2594 & ~w2598) | (~w2594 & w7606) | (~w2598 & w7606);
assign w2774 = ~w2755 & w2773;
assign w2775 = (~w2770 & ~w2755) | (~w2770 & w8410) | (~w2755 & w8410);
assign w2776 = ~w2774 & w2775;
assign w2777 = (~w2616 & ~w2642) | (~w2616 & w8411) | (~w2642 & w8411);
assign w2778 = (~w2660 & ~w2687) | (~w2660 & w8412) | (~w2687 & w8412);
assign w2779 = ~w2777 & ~w2778;
assign w2780 = w2777 & w2778;
assign w2781 = ~w2779 & ~w2780;
assign w2782 = pi03 & ~w2206;
assign w2783 = pi04 & w2032;
assign w2784 = (pi57 & w2782) | (pi57 & w8413) | (w2782 & w8413);
assign w2785 = ~w2782 & w8414;
assign w2786 = ~w2784 & ~w2785;
assign w2787 = (~w2639 & ~w2624) | (~w2639 & w8415) | (~w2624 & w8415);
assign w2788 = ~w2631 & ~w2787;
assign w2789 = ~w2787 & w7607;
assign w2790 = ~w2786 & ~w2788;
assign w2791 = ~w2789 & ~w2790;
assign w2792 = pi10 & w1132;
assign w2793 = pi09 & ~w2419;
assign w2794 = ~w2418 & w2793;
assign w2795 = ~w2792 & ~w2794;
assign w2796 = pi51 & ~w2795;
assign w2797 = ~pi51 & w2795;
assign w2798 = ~w2796 & ~w2797;
assign w2799 = pi06 & w1695;
assign w2800 = (pi55 & ~w1693) | (pi55 & w7608) | (~w1693 & w7608);
assign w2801 = w1694 & w8416;
assign w2802 = ~w2799 & w8417;
assign w2803 = w1695 & w9026;
assign w2804 = ~w2802 & ~w2803;
assign w2805 = ~w2798 & ~w2804;
assign w2806 = w2798 & w2804;
assign w2807 = ~w2805 & ~w2806;
assign w2808 = pi08 & w1393;
assign w2809 = (pi53 & ~w1391) | (pi53 & w8418) | (~w1391 & w8418);
assign w2810 = w1392 & w9027;
assign w2811 = ~w2808 & ~w2809;
assign w2812 = w1393 & w8419;
assign w2813 = (~w2812 & ~w2811) | (~w2812 & w8420) | (~w2811 & w8420);
assign w2814 = w2807 & ~w2813;
assign w2815 = ~w2807 & w2813;
assign w2816 = ~w2814 & ~w2815;
assign w2817 = w2791 & ~w2816;
assign w2818 = ~w2791 & w2816;
assign w2819 = ~w2817 & ~w2818;
assign w2820 = ~w2781 & ~w2819;
assign w2821 = w2781 & w2819;
assign w2822 = ~w2820 & ~w2821;
assign w2823 = ~w2692 & ~w2749;
assign w2824 = ~w2691 & ~w2823;
assign w2825 = ~w2822 & ~w2824;
assign w2826 = w2822 & w2824;
assign w2827 = ~w2825 & ~w2826;
assign w2828 = (~w2684 & ~w2669) | (~w2684 & w8421) | (~w2669 & w8421);
assign w2829 = ~w2676 & ~w2828;
assign w2830 = (~w2743 & ~w2728) | (~w2743 & w8422) | (~w2728 & w8422);
assign w2831 = ~w2735 & ~w2830;
assign w2832 = ~w2829 & ~w2831;
assign w2833 = w2829 & w2831;
assign w2834 = ~w2832 & ~w2833;
assign w2835 = pi16 & w523;
assign w2836 = pi15 & ~w1570;
assign w2837 = ~w1569 & w2836;
assign w2838 = ~w2835 & ~w2837;
assign w2839 = pi45 & ~w2838;
assign w2840 = ~pi45 & w2838;
assign w2841 = ~w2839 & ~w2840;
assign w2842 = pi12 & w909;
assign w2843 = (pi49 & ~w907) | (pi49 & w7609) | (~w907 & w7609);
assign w2844 = w908 & w8423;
assign w2845 = ~w2842 & w8424;
assign w2846 = w909 & w9028;
assign w2847 = ~w2845 & ~w2846;
assign w2848 = ~w2841 & ~w2847;
assign w2849 = w2841 & w2847;
assign w2850 = ~w2848 & ~w2849;
assign w2851 = pi14 & w700;
assign w2852 = (pi47 & ~w698) | (pi47 & w8425) | (~w698 & w8425);
assign w2853 = w699 & w9029;
assign w2854 = ~w2851 & ~w2852;
assign w2855 = w700 & w8426;
assign w2856 = (~w2855 & ~w2854) | (~w2855 & w8427) | (~w2854 & w8427);
assign w2857 = w2850 & ~w2856;
assign w2858 = ~w2850 & w2856;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = w2834 & ~w2859;
assign w2861 = ~w2834 & w2859;
assign w2862 = ~w2860 & ~w2861;
assign w2863 = ~w2719 & w2746;
assign w2864 = ~w2720 & ~w2863;
assign w2865 = ~w2862 & ~w2864;
assign w2866 = w2862 & w2864;
assign w2867 = ~w2865 & ~w2866;
assign w2868 = (~w2707 & ~w2709) | (~w2707 & w7610) | (~w2709 & w7610);
assign w2869 = pi26 & w8;
assign w2870 = (pi35 & ~w6) | (pi35 & w8428) | (~w6 & w8428);
assign w2871 = pi25 & w7;
assign w2872 = ~w2869 & w8429;
assign w2873 = w8 & w9030;
assign w2874 = ~w2872 & ~w2873;
assign w2875 = pi24 & w56;
assign w2876 = (pi37 & ~w54) | (pi37 & w8430) | (~w54 & w8430);
assign w2877 = pi23 & w55;
assign w2878 = ~w2875 & w8431;
assign w2879 = w56 & w9031;
assign w2880 = ~w2878 & ~w2879;
assign w2881 = w2874 & w2880;
assign w2882 = ~w2874 & ~w2880;
assign w2883 = ~w2881 & ~w2882;
assign w2884 = pi28 & pi32;
assign w2885 = pi27 & ~pi32;
assign w2886 = pi33 & ~w2884;
assign w2887 = ~w2885 & w2886;
assign w2888 = ~pi33 & w2884;
assign w2889 = ~w2887 & ~w2888;
assign w2890 = w2883 & ~w2889;
assign w2891 = ~w2883 & w2889;
assign w2892 = ~w2890 & ~w2891;
assign w2893 = ~w2868 & w2892;
assign w2894 = w2868 & ~w2892;
assign w2895 = ~w2893 & ~w2894;
assign w2896 = pi22 & w119;
assign w2897 = pi21 & ~w1634;
assign w2898 = ~w1633 & w2897;
assign w2899 = ~w2896 & ~w2898;
assign w2900 = pi39 & ~w2899;
assign w2901 = ~pi39 & w2899;
assign w2902 = ~w2900 & ~w2901;
assign w2903 = pi20 & w217;
assign w2904 = (pi41 & ~w215) | (pi41 & w8432) | (~w215 & w8432);
assign w2905 = pi19 & w216;
assign w2906 = ~w2903 & w8433;
assign w2907 = w217 & w9032;
assign w2908 = ~w2906 & ~w2907;
assign w2909 = ~w2902 & ~w2908;
assign w2910 = w2902 & w2908;
assign w2911 = ~w2909 & ~w2910;
assign w2912 = pi18 & w355;
assign w2913 = (pi43 & ~w353) | (pi43 & w8434) | (~w353 & w8434);
assign w2914 = pi17 & w354;
assign w2915 = ~w2912 & w8435;
assign w2916 = w355 & w9033;
assign w2917 = ~w2915 & ~w2916;
assign w2918 = w2911 & ~w2917;
assign w2919 = ~w2911 & w2917;
assign w2920 = ~w2918 & ~w2919;
assign w2921 = w2895 & ~w2920;
assign w2922 = ~w2895 & w2920;
assign w2923 = ~w2921 & ~w2922;
assign w2924 = w2867 & ~w2923;
assign w2925 = ~w2867 & w2923;
assign w2926 = ~w2924 & ~w2925;
assign w2927 = ~w2827 & w2926;
assign w2928 = w2827 & ~w2926;
assign w2929 = ~w2927 & ~w2928;
assign w2930 = ~pi59 & ~pi60;
assign w2931 = pi59 & pi60;
assign w2932 = ~w2930 & ~w2931;
assign w2933 = pi00 & w2932;
assign w2934 = pi01 & ~w2588;
assign w2935 = pi02 & w2390;
assign w2936 = (pi59 & w2934) | (pi59 & w8436) | (w2934 & w8436);
assign w2937 = ~w2934 & w8437;
assign w2938 = ~w2936 & ~w2937;
assign w2939 = w2933 & w2938;
assign w2940 = ~w2933 & ~w2938;
assign w2941 = ~w2939 & ~w2940;
assign w2942 = (pi59 & ~w2390) | (pi59 & w8438) | (~w2390 & w8438);
assign w2943 = ~w2589 & w8439;
assign w2944 = ~w2941 & ~w2943;
assign w2945 = w2941 & w2943;
assign w2946 = ~w2944 & ~w2945;
assign w2947 = (~w2605 & ~w2607) | (~w2605 & w8440) | (~w2607 & w8440);
assign w2948 = ~w2946 & w2947;
assign w2949 = w2946 & ~w2947;
assign w2950 = ~w2948 & ~w2949;
assign w2951 = ~w2651 & w2752;
assign w2952 = ~w2652 & ~w2951;
assign w2953 = ~w2951 & w8441;
assign w2954 = (~w2950 & w2951) | (~w2950 & w8442) | (w2951 & w8442);
assign w2955 = ~w2953 & ~w2954;
assign w2956 = w2929 & ~w2955;
assign w2957 = ~w2929 & w2955;
assign w2958 = ~w2956 & ~w2957;
assign w2959 = w2776 & ~w2958;
assign w2960 = ~w2776 & w2958;
assign w2961 = ~w2959 & ~w2960;
assign w2962 = ~w2769 & w2961;
assign w2963 = w2769 & ~w2961;
assign w2964 = ~w2962 & ~w2963;
assign w2965 = ~w2568 & ~w2762;
assign w2966 = (w2761 & w2762) | (w2761 & w8443) | (w2762 & w8443);
assign w2967 = w2569 & w2764;
assign w2968 = ~w2966 & ~w2967;
assign w2969 = ~w2966 & w9080;
assign w2970 = (w2964 & w2969) | (w2964 & w8444) | (w2969 & w8444);
assign w2971 = ~w2969 & w8445;
assign w2972 = ~w2970 & ~w2971;
assign w2973 = ~w2772 & ~w2959;
assign w2974 = (~w2945 & w2947) | (~w2945 & w8446) | (w2947 & w8446);
assign w2975 = w2929 & ~w2954;
assign w2976 = ~w2975 & w7611;
assign w2977 = (~w2974 & w2975) | (~w2974 & w7612) | (w2975 & w7612);
assign w2978 = ~w2976 & ~w2977;
assign w2979 = pi61 & w2930;
assign w2980 = ~pi61 & w2931;
assign w2981 = ~w2979 & ~w2980;
assign w2982 = pi00 & ~w2981;
assign w2983 = pi01 & w2932;
assign w2984 = (pi61 & w2982) | (pi61 & w8447) | (w2982 & w8447);
assign w2985 = ~w2982 & w8448;
assign w2986 = ~w2984 & ~w2985;
assign w2987 = pi02 & ~w2588;
assign w2988 = pi03 & w2390;
assign w2989 = (pi59 & w2987) | (pi59 & w8449) | (w2987 & w8449);
assign w2990 = ~w2987 & w8450;
assign w2991 = ~w2989 & ~w2990;
assign w2992 = w2986 & w2991;
assign w2993 = ~w2986 & ~w2991;
assign w2994 = ~w2992 & ~w2993;
assign w2995 = (pi61 & ~w2932) | (pi61 & w8451) | (~w2932 & w8451);
assign w2996 = (~w2995 & ~w2938) | (~w2995 & w8452) | (~w2938 & w8452);
assign w2997 = ~w2994 & w2996;
assign w2998 = w2994 & ~w2996;
assign w2999 = ~w2997 & ~w2998;
assign w3000 = (~w2780 & ~w2781) | (~w2780 & w8453) | (~w2781 & w8453);
assign w3001 = w2999 & ~w3000;
assign w3002 = ~w2999 & w3000;
assign w3003 = ~w3001 & ~w3002;
assign w3004 = (~w2826 & ~w2827) | (~w2826 & w7613) | (~w2827 & w7613);
assign w3005 = ~w3003 & w3004;
assign w3006 = w3003 & ~w3004;
assign w3007 = ~w3005 & ~w3006;
assign w3008 = (~w2790 & ~w2816) | (~w2790 & w8454) | (~w2816 & w8454);
assign w3009 = (~w2832 & ~w2859) | (~w2832 & w8455) | (~w2859 & w8455);
assign w3010 = w3008 & w3009;
assign w3011 = ~w3008 & ~w3009;
assign w3012 = ~w3010 & ~w3011;
assign w3013 = pi04 & ~w2206;
assign w3014 = pi05 & w2032;
assign w3015 = (pi57 & w3013) | (pi57 & w8456) | (w3013 & w8456);
assign w3016 = ~w3013 & w8457;
assign w3017 = ~w3015 & ~w3016;
assign w3018 = (~w2813 & ~w2798) | (~w2813 & w8458) | (~w2798 & w8458);
assign w3019 = ~w2805 & ~w3018;
assign w3020 = ~w3018 & w7614;
assign w3021 = ~w3017 & ~w3019;
assign w3022 = ~w3020 & ~w3021;
assign w3023 = pi11 & w1132;
assign w3024 = pi10 & ~w2419;
assign w3025 = ~w2418 & w3024;
assign w3026 = ~w3023 & ~w3025;
assign w3027 = pi51 & ~w3026;
assign w3028 = ~pi51 & w3026;
assign w3029 = ~w3027 & ~w3028;
assign w3030 = pi09 & w1393;
assign w3031 = (pi53 & ~w1391) | (pi53 & w8459) | (~w1391 & w8459);
assign w3032 = pi08 & w1392;
assign w3033 = ~w3030 & w8460;
assign w3034 = w1393 & w9034;
assign w3035 = ~w3033 & ~w3034;
assign w3036 = ~w3029 & ~w3035;
assign w3037 = w3029 & w3035;
assign w3038 = ~w3036 & ~w3037;
assign w3039 = pi07 & w1695;
assign w3040 = (pi55 & ~w1693) | (pi55 & w8461) | (~w1693 & w8461);
assign w3041 = pi06 & w1694;
assign w3042 = ~w3039 & w8462;
assign w3043 = w1695 & w9035;
assign w3044 = ~w3042 & ~w3043;
assign w3045 = w3038 & ~w3044;
assign w3046 = ~w3038 & w3044;
assign w3047 = ~w3045 & ~w3046;
assign w3048 = w3022 & ~w3047;
assign w3049 = ~w3022 & w3047;
assign w3050 = ~w3048 & ~w3049;
assign w3051 = ~w3012 & w3050;
assign w3052 = w3012 & ~w3050;
assign w3053 = ~w3051 & ~w3052;
assign w3054 = ~w2866 & ~w2923;
assign w3055 = ~w2865 & ~w3054;
assign w3056 = w3053 & ~w3055;
assign w3057 = ~w3053 & w3055;
assign w3058 = ~w3056 & ~w3057;
assign w3059 = (~w2917 & ~w2902) | (~w2917 & w8463) | (~w2902 & w8463);
assign w3060 = ~w2909 & ~w3059;
assign w3061 = (~w2856 & ~w2841) | (~w2856 & w8464) | (~w2841 & w8464);
assign w3062 = ~w2848 & ~w3061;
assign w3063 = ~w3060 & ~w3062;
assign w3064 = w3060 & w3062;
assign w3065 = ~w3063 & ~w3064;
assign w3066 = pi17 & w523;
assign w3067 = pi16 & ~w1570;
assign w3068 = ~w1569 & w3067;
assign w3069 = ~w3066 & ~w3068;
assign w3070 = pi45 & ~w3069;
assign w3071 = ~pi45 & w3069;
assign w3072 = ~w3070 & ~w3071;
assign w3073 = pi13 & w909;
assign w3074 = (pi49 & ~w907) | (pi49 & w8465) | (~w907 & w8465);
assign w3075 = pi12 & w908;
assign w3076 = ~w3073 & w8466;
assign w3077 = w909 & w9036;
assign w3078 = ~w3076 & ~w3077;
assign w3079 = ~w3072 & ~w3078;
assign w3080 = w3072 & w3078;
assign w3081 = ~w3079 & ~w3080;
assign w3082 = pi15 & w700;
assign w3083 = (pi47 & ~w698) | (pi47 & w8467) | (~w698 & w8467);
assign w3084 = pi14 & w699;
assign w3085 = ~w3082 & w8468;
assign w3086 = w700 & w9037;
assign w3087 = ~w3085 & ~w3086;
assign w3088 = w3081 & ~w3087;
assign w3089 = ~w3081 & w3087;
assign w3090 = ~w3088 & ~w3089;
assign w3091 = w3065 & ~w3090;
assign w3092 = ~w3065 & w3090;
assign w3093 = ~w3091 & ~w3092;
assign w3094 = ~w2893 & w2920;
assign w3095 = ~w2894 & ~w3094;
assign w3096 = ~w3093 & ~w3095;
assign w3097 = w3093 & w3095;
assign w3098 = ~w3096 & ~w3097;
assign w3099 = (~w2881 & ~w2883) | (~w2881 & w7615) | (~w2883 & w7615);
assign w3100 = pi25 & w56;
assign w3101 = (pi37 & ~w54) | (pi37 & w8469) | (~w54 & w8469);
assign w3102 = pi24 & w55;
assign w3103 = ~w3100 & w8470;
assign w3104 = w56 & w9038;
assign w3105 = ~w3103 & ~w3104;
assign w3106 = pi27 & w8;
assign w3107 = (pi35 & ~w6) | (pi35 & w8471) | (~w6 & w8471);
assign w3108 = pi26 & w7;
assign w3109 = ~w3106 & w8472;
assign w3110 = w8 & w9039;
assign w3111 = ~w3109 & ~w3110;
assign w3112 = w3105 & w3111;
assign w3113 = ~w3105 & ~w3111;
assign w3114 = ~w3112 & ~w3113;
assign w3115 = pi29 & pi32;
assign w3116 = pi28 & ~pi32;
assign w3117 = pi33 & ~w3115;
assign w3118 = ~w3116 & w3117;
assign w3119 = ~pi33 & w3115;
assign w3120 = ~w3118 & ~w3119;
assign w3121 = w3114 & ~w3120;
assign w3122 = ~w3114 & w3120;
assign w3123 = ~w3121 & ~w3122;
assign w3124 = ~w3099 & w3123;
assign w3125 = w3099 & ~w3123;
assign w3126 = ~w3124 & ~w3125;
assign w3127 = pi23 & w119;
assign w3128 = pi22 & ~w1634;
assign w3129 = ~w1633 & w3128;
assign w3130 = ~w3127 & ~w3129;
assign w3131 = pi39 & ~w3130;
assign w3132 = ~pi39 & w3130;
assign w3133 = ~w3131 & ~w3132;
assign w3134 = pi21 & w217;
assign w3135 = (pi41 & ~w215) | (pi41 & w8473) | (~w215 & w8473);
assign w3136 = pi20 & w216;
assign w3137 = ~w3134 & w8474;
assign w3138 = w217 & w9040;
assign w3139 = ~w3137 & ~w3138;
assign w3140 = ~w3133 & ~w3139;
assign w3141 = w3133 & w3139;
assign w3142 = ~w3140 & ~w3141;
assign w3143 = pi19 & w355;
assign w3144 = (pi43 & ~w353) | (pi43 & w8475) | (~w353 & w8475);
assign w3145 = pi18 & w354;
assign w3146 = ~w3143 & w8476;
assign w3147 = w355 & w9041;
assign w3148 = ~w3146 & ~w3147;
assign w3149 = w3142 & ~w3148;
assign w3150 = ~w3142 & w3148;
assign w3151 = ~w3149 & ~w3150;
assign w3152 = w3126 & ~w3151;
assign w3153 = ~w3126 & w3151;
assign w3154 = ~w3152 & ~w3153;
assign w3155 = w3098 & ~w3154;
assign w3156 = ~w3098 & w3154;
assign w3157 = ~w3155 & ~w3156;
assign w3158 = w3058 & ~w3157;
assign w3159 = ~w3058 & w3157;
assign w3160 = ~w3158 & ~w3159;
assign w3161 = w3007 & ~w3160;
assign w3162 = ~w3007 & w3160;
assign w3163 = ~w3161 & ~w3162;
assign w3164 = w2978 & ~w3163;
assign w3165 = ~w2978 & w3163;
assign w3166 = ~w3164 & ~w3165;
assign w3167 = ~w2973 & w3166;
assign w3168 = w2973 & ~w3166;
assign w3169 = ~w3167 & ~w3168;
assign w3170 = w2764 & w8477;
assign w3171 = (~w2962 & w2965) | (~w2962 & w7616) | (w2965 & w7616);
assign w3172 = ~w3170 & w3171;
assign w3173 = (~w2963 & w3170) | (~w2963 & w7617) | (w3170 & w7617);
assign w3174 = w2371 & w2964;
assign w3175 = w2967 & w3174;
assign w3176 = w3169 & w9081;
assign w3177 = ~w3173 & w9082;
assign w3178 = ~w3176 & ~w3177;
assign w3179 = ~w3005 & w3160;
assign w3180 = w3001 & w3179;
assign w3181 = (~w3001 & w3004) | (~w3001 & w7888) | (w3004 & w7888);
assign w3182 = ~w3179 & w3181;
assign w3183 = ~w3180 & ~w3182;
assign w3184 = ~pi61 & ~pi62;
assign w3185 = pi61 & pi62;
assign w3186 = ~w3184 & ~w3185;
assign w3187 = (pi63 & ~w3186) | (pi63 & w8479) | (~w3186 & w8479);
assign w3188 = w3186 & w8480;
assign w3189 = ~w3187 & ~w3188;
assign w3190 = pi01 & ~w2981;
assign w3191 = pi02 & w2932;
assign w3192 = (pi61 & w3190) | (pi61 & w8481) | (w3190 & w8481);
assign w3193 = ~w3190 & w8482;
assign w3194 = ~w3192 & ~w3193;
assign w3195 = w3189 & ~w3194;
assign w3196 = ~w3189 & w3194;
assign w3197 = ~w3195 & ~w3196;
assign w3198 = pi03 & ~w2588;
assign w3199 = pi04 & w2390;
assign w3200 = (pi59 & w3198) | (pi59 & w8483) | (w3198 & w8483);
assign w3201 = ~w3198 & w8484;
assign w3202 = ~w3200 & ~w3201;
assign w3203 = w3197 & ~w3202;
assign w3204 = ~w3197 & w3202;
assign w3205 = ~w3203 & ~w3204;
assign w3206 = pi63 & w2992;
assign w3207 = ~pi63 & ~w2992;
assign w3208 = ~w3206 & ~w3207;
assign w3209 = ~w3205 & w3208;
assign w3210 = w3205 & ~w3208;
assign w3211 = ~w3209 & ~w3210;
assign w3212 = w2998 & w3211;
assign w3213 = ~w2998 & ~w3211;
assign w3214 = ~w3212 & ~w3213;
assign w3215 = (~w3011 & ~w3012) | (~w3011 & w8485) | (~w3012 & w8485);
assign w3216 = w3214 & w3215;
assign w3217 = ~w3214 & ~w3215;
assign w3218 = ~w3216 & ~w3217;
assign w3219 = ~w3057 & w3157;
assign w3220 = ~w3056 & ~w3219;
assign w3221 = (~w3218 & w3219) | (~w3218 & w8486) | (w3219 & w8486);
assign w3222 = ~w3219 & w8487;
assign w3223 = ~w3221 & ~w3222;
assign w3224 = (~w3021 & ~w3047) | (~w3021 & w8488) | (~w3047 & w8488);
assign w3225 = (~w3063 & ~w3090) | (~w3063 & w8489) | (~w3090 & w8489);
assign w3226 = w3224 & w3225;
assign w3227 = ~w3224 & ~w3225;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = pi05 & ~w2206;
assign w3230 = pi06 & w2032;
assign w3231 = (pi57 & w3229) | (pi57 & w8490) | (w3229 & w8490);
assign w3232 = ~w3229 & w8491;
assign w3233 = ~w3231 & ~w3232;
assign w3234 = (~w3044 & ~w3029) | (~w3044 & w8492) | (~w3029 & w8492);
assign w3235 = ~w3036 & ~w3234;
assign w3236 = ~w3233 & ~w3235;
assign w3237 = ~w3234 & w7618;
assign w3238 = ~w3236 & ~w3237;
assign w3239 = pi12 & w1132;
assign w3240 = pi11 & ~w2419;
assign w3241 = ~w2418 & w3240;
assign w3242 = ~w3239 & ~w3241;
assign w3243 = pi51 & ~w3242;
assign w3244 = ~pi51 & w3242;
assign w3245 = ~w3243 & ~w3244;
assign w3246 = pi10 & w1393;
assign w3247 = (pi53 & ~w1391) | (pi53 & w8493) | (~w1391 & w8493);
assign w3248 = pi09 & w1392;
assign w3249 = ~w3246 & w8494;
assign w3250 = w1393 & w9042;
assign w3251 = ~w3249 & ~w3250;
assign w3252 = ~w3245 & ~w3251;
assign w3253 = w3245 & w3251;
assign w3254 = ~w3252 & ~w3253;
assign w3255 = pi08 & w1695;
assign w3256 = (pi55 & ~w1693) | (pi55 & w8495) | (~w1693 & w8495);
assign w3257 = pi07 & w1694;
assign w3258 = ~w3255 & w8496;
assign w3259 = w1695 & w9043;
assign w3260 = ~w3258 & ~w3259;
assign w3261 = w3254 & ~w3260;
assign w3262 = ~w3254 & w3260;
assign w3263 = ~w3261 & ~w3262;
assign w3264 = w3238 & ~w3263;
assign w3265 = ~w3238 & w3263;
assign w3266 = ~w3264 & ~w3265;
assign w3267 = ~w3228 & w3266;
assign w3268 = w3228 & ~w3266;
assign w3269 = ~w3267 & ~w3268;
assign w3270 = ~w3097 & ~w3154;
assign w3271 = ~w3096 & ~w3270;
assign w3272 = w3269 & ~w3271;
assign w3273 = ~w3269 & w3271;
assign w3274 = ~w3272 & ~w3273;
assign w3275 = (~w3087 & ~w3072) | (~w3087 & w8497) | (~w3072 & w8497);
assign w3276 = ~w3079 & ~w3275;
assign w3277 = (~w3148 & ~w3133) | (~w3148 & w8498) | (~w3133 & w8498);
assign w3278 = ~w3140 & ~w3277;
assign w3279 = w3276 & w3278;
assign w3280 = ~w3276 & ~w3278;
assign w3281 = ~w3279 & ~w3280;
assign w3282 = pi18 & w523;
assign w3283 = pi17 & ~w1570;
assign w3284 = ~w1569 & w3283;
assign w3285 = ~w3282 & ~w3284;
assign w3286 = pi45 & ~w3285;
assign w3287 = ~pi45 & w3285;
assign w3288 = ~w3286 & ~w3287;
assign w3289 = pi14 & w909;
assign w3290 = (pi49 & ~w907) | (pi49 & w8499) | (~w907 & w8499);
assign w3291 = pi13 & w908;
assign w3292 = ~w3289 & w8500;
assign w3293 = w909 & w9044;
assign w3294 = ~w3292 & ~w3293;
assign w3295 = ~w3288 & ~w3294;
assign w3296 = w3288 & w3294;
assign w3297 = ~w3295 & ~w3296;
assign w3298 = pi16 & w700;
assign w3299 = (pi47 & ~w698) | (pi47 & w8501) | (~w698 & w8501);
assign w3300 = pi15 & w699;
assign w3301 = ~w3298 & w8502;
assign w3302 = w700 & w9045;
assign w3303 = ~w3301 & ~w3302;
assign w3304 = w3297 & ~w3303;
assign w3305 = ~w3297 & w3303;
assign w3306 = ~w3304 & ~w3305;
assign w3307 = w3281 & w3306;
assign w3308 = ~w3281 & ~w3306;
assign w3309 = ~w3307 & ~w3308;
assign w3310 = ~w3124 & w3151;
assign w3311 = ~w3125 & ~w3310;
assign w3312 = ~w3309 & w3311;
assign w3313 = w3309 & ~w3311;
assign w3314 = ~w3312 & ~w3313;
assign w3315 = (~w3112 & ~w3114) | (~w3112 & w7619) | (~w3114 & w7619);
assign w3316 = pi26 & w56;
assign w3317 = (pi37 & ~w54) | (pi37 & w8503) | (~w54 & w8503);
assign w3318 = pi25 & w55;
assign w3319 = ~w3316 & w8504;
assign w3320 = w56 & w9046;
assign w3321 = ~w3319 & ~w3320;
assign w3322 = pi28 & w8;
assign w3323 = (pi35 & ~w6) | (pi35 & w8505) | (~w6 & w8505);
assign w3324 = pi27 & w7;
assign w3325 = ~w3322 & w8506;
assign w3326 = w8 & w9047;
assign w3327 = ~w3325 & ~w3326;
assign w3328 = w3321 & w3327;
assign w3329 = ~w3321 & ~w3327;
assign w3330 = ~w3328 & ~w3329;
assign w3331 = pi30 & pi32;
assign w3332 = pi29 & ~pi32;
assign w3333 = pi33 & ~w3331;
assign w3334 = ~w3332 & w3333;
assign w3335 = ~pi33 & w3331;
assign w3336 = ~w3334 & ~w3335;
assign w3337 = w3330 & ~w3336;
assign w3338 = ~w3330 & w3336;
assign w3339 = ~w3337 & ~w3338;
assign w3340 = ~w3315 & w3339;
assign w3341 = w3315 & ~w3339;
assign w3342 = ~w3340 & ~w3341;
assign w3343 = pi24 & w119;
assign w3344 = pi23 & ~w1634;
assign w3345 = ~w1633 & w3344;
assign w3346 = ~w3343 & ~w3345;
assign w3347 = pi39 & ~w3346;
assign w3348 = ~pi39 & w3346;
assign w3349 = ~w3347 & ~w3348;
assign w3350 = pi22 & w217;
assign w3351 = (pi41 & ~w215) | (pi41 & w8507) | (~w215 & w8507);
assign w3352 = pi21 & w216;
assign w3353 = ~w3350 & w8508;
assign w3354 = w217 & w9048;
assign w3355 = ~w3353 & ~w3354;
assign w3356 = ~w3349 & ~w3355;
assign w3357 = w3349 & w3355;
assign w3358 = ~w3356 & ~w3357;
assign w3359 = pi20 & w355;
assign w3360 = (pi43 & ~w353) | (pi43 & w8509) | (~w353 & w8509);
assign w3361 = pi19 & w354;
assign w3362 = ~w3359 & w8510;
assign w3363 = w355 & w9049;
assign w3364 = ~w3362 & ~w3363;
assign w3365 = w3358 & ~w3364;
assign w3366 = ~w3358 & w3364;
assign w3367 = ~w3365 & ~w3366;
assign w3368 = w3342 & ~w3367;
assign w3369 = ~w3342 & w3367;
assign w3370 = ~w3368 & ~w3369;
assign w3371 = w3314 & ~w3370;
assign w3372 = ~w3314 & w3370;
assign w3373 = ~w3371 & ~w3372;
assign w3374 = w3274 & ~w3373;
assign w3375 = ~w3274 & w3373;
assign w3376 = ~w3374 & ~w3375;
assign w3377 = w3223 & ~w3376;
assign w3378 = ~w3223 & w3376;
assign w3379 = ~w3377 & ~w3378;
assign w3380 = ~w3183 & w3379;
assign w3381 = w3183 & ~w3379;
assign w3382 = ~w3380 & ~w3381;
assign w3383 = ~w2977 & ~w3164;
assign w3384 = w3382 & ~w3383;
assign w3385 = ~w3382 & w3383;
assign w3386 = ~w3384 & ~w3385;
assign w3387 = ~w3176 & w8511;
assign w3388 = (w3386 & w3176) | (w3386 & w8512) | (w3176 & w8512);
assign w3389 = ~w3387 & ~w3388;
assign w3390 = (~w3180 & ~w3183) | (~w3180 & w8513) | (~w3183 & w8513);
assign w3391 = ~w3212 & ~w3216;
assign w3392 = ~w3221 & w3376;
assign w3393 = (~w3391 & w3392) | (~w3391 & w7620) | (w3392 & w7620);
assign w3394 = ~w3392 & w7621;
assign w3395 = ~w3393 & ~w3394;
assign w3396 = (~w3195 & ~w3197) | (~w3195 & w8514) | (~w3197 & w8514);
assign w3397 = pi04 & ~w2588;
assign w3398 = pi05 & w2390;
assign w3399 = (pi59 & w3397) | (pi59 & w8515) | (w3397 & w8515);
assign w3400 = ~w3397 & w8516;
assign w3401 = ~w3399 & ~w3400;
assign w3402 = pi63 & w3184;
assign w3403 = ~pi63 & w3185;
assign w3404 = ~w3402 & ~w3403;
assign w3405 = pi00 & ~w3404;
assign w3406 = pi01 & w3186;
assign w3407 = (pi63 & w3405) | (pi63 & w8517) | (w3405 & w8517);
assign w3408 = ~w3405 & w8518;
assign w3409 = ~w3407 & ~w3408;
assign w3410 = pi02 & ~w2981;
assign w3411 = pi03 & w2932;
assign w3412 = (pi61 & w3410) | (pi61 & w8519) | (w3410 & w8519);
assign w3413 = ~w3410 & w8520;
assign w3414 = ~w3412 & ~w3413;
assign w3415 = w3409 & w3414;
assign w3416 = ~w3409 & ~w3414;
assign w3417 = ~w3415 & ~w3416;
assign w3418 = w3401 & w3417;
assign w3419 = ~w3401 & ~w3417;
assign w3420 = ~w3418 & ~w3419;
assign w3421 = w3396 & w3420;
assign w3422 = ~w3396 & ~w3420;
assign w3423 = ~w3421 & ~w3422;
assign w3424 = (~w3206 & w3205) | (~w3206 & w8521) | (w3205 & w8521);
assign w3425 = w3423 & ~w3424;
assign w3426 = ~w3423 & w3424;
assign w3427 = ~w3425 & ~w3426;
assign w3428 = (~w3227 & ~w3228) | (~w3227 & w8522) | (~w3228 & w8522);
assign w3429 = w3427 & w3428;
assign w3430 = ~w3427 & ~w3428;
assign w3431 = ~w3429 & ~w3430;
assign w3432 = ~w3273 & w3373;
assign w3433 = ~w3272 & ~w3432;
assign w3434 = (~w3431 & w3432) | (~w3431 & w8523) | (w3432 & w8523);
assign w3435 = ~w3432 & w8524;
assign w3436 = ~w3434 & ~w3435;
assign w3437 = (~w3279 & w3306) | (~w3279 & w8525) | (w3306 & w8525);
assign w3438 = (~w3236 & ~w3263) | (~w3236 & w8526) | (~w3263 & w8526);
assign w3439 = w3437 & ~w3438;
assign w3440 = ~w3437 & w3438;
assign w3441 = ~w3439 & ~w3440;
assign w3442 = pi06 & ~w2206;
assign w3443 = pi07 & w2032;
assign w3444 = (pi57 & w3442) | (pi57 & w8527) | (w3442 & w8527);
assign w3445 = ~w3442 & w8528;
assign w3446 = ~w3444 & ~w3445;
assign w3447 = (~w3260 & ~w3245) | (~w3260 & w8529) | (~w3245 & w8529);
assign w3448 = ~w3252 & ~w3447;
assign w3449 = ~w3447 & w7622;
assign w3450 = ~w3446 & ~w3448;
assign w3451 = ~w3449 & ~w3450;
assign w3452 = pi13 & w1132;
assign w3453 = pi12 & ~w2419;
assign w3454 = ~w2418 & w3453;
assign w3455 = ~w3452 & ~w3454;
assign w3456 = pi51 & ~w3455;
assign w3457 = ~pi51 & w3455;
assign w3458 = ~w3456 & ~w3457;
assign w3459 = pi11 & w1393;
assign w3460 = (pi53 & ~w1391) | (pi53 & w8530) | (~w1391 & w8530);
assign w3461 = pi10 & w1392;
assign w3462 = ~w3459 & w8531;
assign w3463 = pi53 & w3459;
assign w3464 = ~w3462 & ~w3463;
assign w3465 = ~w3458 & ~w3464;
assign w3466 = w3458 & w3464;
assign w3467 = ~w3465 & ~w3466;
assign w3468 = pi09 & w1695;
assign w3469 = (pi55 & ~w1693) | (pi55 & w8532) | (~w1693 & w8532);
assign w3470 = pi08 & w1694;
assign w3471 = ~w3468 & w8533;
assign w3472 = pi55 & w3468;
assign w3473 = ~w3471 & ~w3472;
assign w3474 = w3467 & ~w3473;
assign w3475 = ~w3467 & w3473;
assign w3476 = ~w3474 & ~w3475;
assign w3477 = w3451 & ~w3476;
assign w3478 = ~w3451 & w3476;
assign w3479 = ~w3477 & ~w3478;
assign w3480 = ~w3441 & w3479;
assign w3481 = w3441 & ~w3479;
assign w3482 = ~w3480 & ~w3481;
assign w3483 = ~w3312 & ~w3370;
assign w3484 = ~w3313 & ~w3483;
assign w3485 = ~w3482 & w3484;
assign w3486 = w3482 & ~w3484;
assign w3487 = ~w3485 & ~w3486;
assign w3488 = (~w3303 & ~w3288) | (~w3303 & w8534) | (~w3288 & w8534);
assign w3489 = ~w3295 & ~w3488;
assign w3490 = (~w3364 & ~w3349) | (~w3364 & w8535) | (~w3349 & w8535);
assign w3491 = ~w3356 & ~w3490;
assign w3492 = ~w3489 & ~w3491;
assign w3493 = w3489 & w3491;
assign w3494 = ~w3492 & ~w3493;
assign w3495 = pi19 & w523;
assign w3496 = pi18 & ~w1570;
assign w3497 = ~w1569 & w3496;
assign w3498 = ~w3495 & ~w3497;
assign w3499 = pi45 & ~w3498;
assign w3500 = ~pi45 & w3498;
assign w3501 = ~w3499 & ~w3500;
assign w3502 = pi17 & w700;
assign w3503 = (pi47 & ~w698) | (pi47 & w8536) | (~w698 & w8536);
assign w3504 = pi16 & w699;
assign w3505 = ~w3502 & w8537;
assign w3506 = pi47 & w3502;
assign w3507 = ~w3505 & ~w3506;
assign w3508 = ~w3501 & ~w3507;
assign w3509 = w3501 & w3507;
assign w3510 = ~w3508 & ~w3509;
assign w3511 = pi15 & w909;
assign w3512 = (pi49 & ~w907) | (pi49 & w8538) | (~w907 & w8538);
assign w3513 = pi14 & w908;
assign w3514 = ~w3511 & w8539;
assign w3515 = pi49 & w3511;
assign w3516 = ~w3514 & ~w3515;
assign w3517 = w3510 & ~w3516;
assign w3518 = ~w3510 & w3516;
assign w3519 = ~w3517 & ~w3518;
assign w3520 = w3494 & ~w3519;
assign w3521 = ~w3494 & w3519;
assign w3522 = ~w3520 & ~w3521;
assign w3523 = ~w3340 & w3367;
assign w3524 = ~w3341 & ~w3523;
assign w3525 = ~w3522 & ~w3524;
assign w3526 = w3522 & w3524;
assign w3527 = ~w3525 & ~w3526;
assign w3528 = (~w3328 & ~w3330) | (~w3328 & w7623) | (~w3330 & w7623);
assign w3529 = pi31 & pi32;
assign w3530 = ~pi33 & w3529;
assign w3531 = pi30 & ~pi32;
assign w3532 = pi33 & ~w3529;
assign w3533 = ~w3531 & w3532;
assign w3534 = ~w3530 & ~w3533;
assign w3535 = pi29 & w8;
assign w3536 = (pi35 & ~w6) | (pi35 & w8540) | (~w6 & w8540);
assign w3537 = pi28 & w7;
assign w3538 = ~w3535 & w8541;
assign w3539 = w8 & w9050;
assign w3540 = ~w3538 & ~w3539;
assign w3541 = pi27 & w56;
assign w3542 = (pi37 & ~w54) | (pi37 & w8542) | (~w54 & w8542);
assign w3543 = pi26 & w55;
assign w3544 = ~w3541 & w8543;
assign w3545 = w56 & w9051;
assign w3546 = ~w3544 & ~w3545;
assign w3547 = w3540 & w3546;
assign w3548 = ~w3540 & ~w3546;
assign w3549 = ~w3547 & ~w3548;
assign w3550 = ~w3534 & w3549;
assign w3551 = w3534 & ~w3549;
assign w3552 = ~w3550 & ~w3551;
assign w3553 = ~w3528 & w3552;
assign w3554 = w3528 & ~w3552;
assign w3555 = ~w3553 & ~w3554;
assign w3556 = pi25 & w119;
assign w3557 = pi24 & ~w1634;
assign w3558 = ~w1633 & w3557;
assign w3559 = ~w3556 & ~w3558;
assign w3560 = pi39 & ~w3559;
assign w3561 = ~pi39 & w3559;
assign w3562 = ~w3560 & ~w3561;
assign w3563 = pi23 & w217;
assign w3564 = (pi41 & ~w215) | (pi41 & w8544) | (~w215 & w8544);
assign w3565 = pi22 & w216;
assign w3566 = ~w3563 & w8545;
assign w3567 = pi41 & w3563;
assign w3568 = ~w3566 & ~w3567;
assign w3569 = ~w3562 & ~w3568;
assign w3570 = w3562 & w3568;
assign w3571 = ~w3569 & ~w3570;
assign w3572 = pi21 & w355;
assign w3573 = (pi43 & ~w353) | (pi43 & w8546) | (~w353 & w8546);
assign w3574 = pi20 & w354;
assign w3575 = ~w3572 & w8547;
assign w3576 = pi43 & w3572;
assign w3577 = ~w3575 & ~w3576;
assign w3578 = w3571 & ~w3577;
assign w3579 = ~w3571 & w3577;
assign w3580 = ~w3578 & ~w3579;
assign w3581 = w3555 & ~w3580;
assign w3582 = ~w3555 & w3580;
assign w3583 = ~w3581 & ~w3582;
assign w3584 = w3527 & ~w3583;
assign w3585 = ~w3527 & w3583;
assign w3586 = ~w3584 & ~w3585;
assign w3587 = w3487 & w3586;
assign w3588 = ~w3487 & ~w3586;
assign w3589 = ~w3587 & ~w3588;
assign w3590 = w3436 & ~w3589;
assign w3591 = ~w3436 & w3589;
assign w3592 = ~w3590 & ~w3591;
assign w3593 = w3395 & w3592;
assign w3594 = ~w3395 & ~w3592;
assign w3595 = ~w3593 & ~w3594;
assign w3596 = w3390 & ~w3595;
assign w3597 = ~w3390 & w3595;
assign w3598 = ~w3596 & ~w3597;
assign w3599 = ~w3168 & ~w3385;
assign w3600 = ~w3384 & ~w3599;
assign w3601 = w3175 & w7889;
assign w3602 = ~w2380 & w3601;
assign w3603 = ~w3167 & ~w3384;
assign w3604 = ~w3385 & ~w3603;
assign w3605 = w3169 & w3386;
assign w3606 = ~w2963 & w3605;
assign w3607 = (~w3604 & w3172) | (~w3604 & w7624) | (w3172 & w7624);
assign w3608 = (w3598 & w3602) | (w3598 & w8548) | (w3602 & w8548);
assign w3609 = ~w3602 & w8549;
assign w3610 = ~w3608 & ~w3609;
assign w3611 = ~w3599 & w8550;
assign w3612 = w3175 & w8551;
assign w3613 = ~w2380 & w3612;
assign w3614 = w2962 & w3605;
assign w3615 = (~w3597 & w3603) | (~w3597 & w7890) | (w3603 & w7890);
assign w3616 = ~w3614 & w3615;
assign w3617 = ~w3173 & w3616;
assign w3618 = (~w3611 & w3173) | (~w3611 & w8552) | (w3173 & w8552);
assign w3619 = ~w3613 & ~w3618;
assign w3620 = (~w3393 & ~w3395) | (~w3393 & w8553) | (~w3395 & w8553);
assign w3621 = ~w3425 & ~w3429;
assign w3622 = ~w3435 & w3589;
assign w3623 = (w3621 & w3622) | (w3621 & w7625) | (w3622 & w7625);
assign w3624 = ~w3622 & w7626;
assign w3625 = ~w3623 & ~w3624;
assign w3626 = (~w3415 & ~w3417) | (~w3415 & w8554) | (~w3417 & w8554);
assign w3627 = pi05 & ~w2588;
assign w3628 = pi06 & w2390;
assign w3629 = (pi59 & w3627) | (pi59 & w8555) | (w3627 & w8555);
assign w3630 = ~w3627 & w8556;
assign w3631 = ~w3629 & ~w3630;
assign w3632 = pi01 & ~w3404;
assign w3633 = pi02 & w3186;
assign w3634 = (pi63 & w3632) | (pi63 & w8557) | (w3632 & w8557);
assign w3635 = ~w3632 & w8558;
assign w3636 = ~w3634 & ~w3635;
assign w3637 = pi03 & ~w2981;
assign w3638 = pi04 & w2932;
assign w3639 = (pi61 & w3637) | (pi61 & w8559) | (w3637 & w8559);
assign w3640 = ~w3637 & w8560;
assign w3641 = ~w3639 & ~w3640;
assign w3642 = w3636 & w3641;
assign w3643 = ~w3636 & ~w3641;
assign w3644 = ~w3642 & ~w3643;
assign w3645 = w3631 & w3644;
assign w3646 = ~w3631 & ~w3644;
assign w3647 = ~w3645 & ~w3646;
assign w3648 = ~w3626 & w3647;
assign w3649 = w3626 & ~w3647;
assign w3650 = ~w3648 & ~w3649;
assign w3651 = w3421 & ~w3650;
assign w3652 = ~w3421 & w3650;
assign w3653 = ~w3651 & ~w3652;
assign w3654 = (~w3439 & ~w3441) | (~w3439 & w8561) | (~w3441 & w8561);
assign w3655 = ~w3653 & ~w3654;
assign w3656 = w3653 & w3654;
assign w3657 = ~w3655 & ~w3656;
assign w3658 = ~w3486 & ~w3586;
assign w3659 = ~w3485 & ~w3658;
assign w3660 = (w3657 & w3658) | (w3657 & w8562) | (w3658 & w8562);
assign w3661 = ~w3658 & w8563;
assign w3662 = ~w3660 & ~w3661;
assign w3663 = (~w3492 & ~w3519) | (~w3492 & w8564) | (~w3519 & w8564);
assign w3664 = (~w3450 & ~w3476) | (~w3450 & w8565) | (~w3476 & w8565);
assign w3665 = ~w3663 & ~w3664;
assign w3666 = w3663 & w3664;
assign w3667 = ~w3665 & ~w3666;
assign w3668 = pi07 & ~w2206;
assign w3669 = pi08 & w2032;
assign w3670 = (pi57 & w3668) | (pi57 & w8566) | (w3668 & w8566);
assign w3671 = ~w3668 & w8567;
assign w3672 = ~w3670 & ~w3671;
assign w3673 = (~w3473 & ~w3458) | (~w3473 & w8568) | (~w3458 & w8568);
assign w3674 = ~w3465 & ~w3673;
assign w3675 = ~w3672 & ~w3674;
assign w3676 = ~w3673 & w7627;
assign w3677 = ~w3675 & ~w3676;
assign w3678 = pi14 & w1132;
assign w3679 = pi13 & ~w2419;
assign w3680 = ~w2418 & w3679;
assign w3681 = ~w3678 & ~w3680;
assign w3682 = pi51 & ~w3681;
assign w3683 = ~pi51 & w3681;
assign w3684 = ~w3682 & ~w3683;
assign w3685 = pi12 & w1393;
assign w3686 = (pi53 & ~w1391) | (pi53 & w8569) | (~w1391 & w8569);
assign w3687 = pi11 & w1392;
assign w3688 = ~w3685 & w8570;
assign w3689 = pi53 & w3685;
assign w3690 = ~w3688 & ~w3689;
assign w3691 = ~w3684 & ~w3690;
assign w3692 = w3684 & w3690;
assign w3693 = ~w3691 & ~w3692;
assign w3694 = pi10 & w1695;
assign w3695 = (pi55 & ~w1693) | (pi55 & w8571) | (~w1693 & w8571);
assign w3696 = pi09 & w1694;
assign w3697 = ~w3694 & w8572;
assign w3698 = pi55 & w3694;
assign w3699 = ~w3697 & ~w3698;
assign w3700 = w3693 & ~w3699;
assign w3701 = ~w3693 & w3699;
assign w3702 = ~w3700 & ~w3701;
assign w3703 = w3677 & ~w3702;
assign w3704 = ~w3677 & w3702;
assign w3705 = ~w3703 & ~w3704;
assign w3706 = ~w3667 & ~w3705;
assign w3707 = w3667 & w3705;
assign w3708 = ~w3706 & ~w3707;
assign w3709 = ~w3526 & ~w3583;
assign w3710 = ~w3525 & ~w3709;
assign w3711 = ~w3708 & ~w3710;
assign w3712 = w3708 & w3710;
assign w3713 = ~w3711 & ~w3712;
assign w3714 = (~w3516 & ~w3501) | (~w3516 & w8573) | (~w3501 & w8573);
assign w3715 = ~w3508 & ~w3714;
assign w3716 = (~w3577 & ~w3562) | (~w3577 & w8574) | (~w3562 & w8574);
assign w3717 = ~w3569 & ~w3716;
assign w3718 = ~w3715 & ~w3717;
assign w3719 = w3715 & w3717;
assign w3720 = ~w3718 & ~w3719;
assign w3721 = pi20 & w523;
assign w3722 = pi19 & ~w1570;
assign w3723 = ~w1569 & w3722;
assign w3724 = ~w3721 & ~w3723;
assign w3725 = pi45 & ~w3724;
assign w3726 = ~pi45 & w3724;
assign w3727 = ~w3725 & ~w3726;
assign w3728 = pi18 & w700;
assign w3729 = (pi47 & ~w698) | (pi47 & w8575) | (~w698 & w8575);
assign w3730 = pi17 & w699;
assign w3731 = ~w3728 & w8576;
assign w3732 = pi47 & w3728;
assign w3733 = ~w3731 & ~w3732;
assign w3734 = ~w3727 & ~w3733;
assign w3735 = w3727 & w3733;
assign w3736 = ~w3734 & ~w3735;
assign w3737 = pi16 & w909;
assign w3738 = (pi49 & ~w907) | (pi49 & w8577) | (~w907 & w8577);
assign w3739 = pi15 & w908;
assign w3740 = ~w3737 & w8578;
assign w3741 = pi49 & w3737;
assign w3742 = ~w3740 & ~w3741;
assign w3743 = w3736 & ~w3742;
assign w3744 = ~w3736 & w3742;
assign w3745 = ~w3743 & ~w3744;
assign w3746 = w3720 & ~w3745;
assign w3747 = ~w3720 & w3745;
assign w3748 = ~w3746 & ~w3747;
assign w3749 = ~w3553 & w3580;
assign w3750 = ~w3554 & ~w3749;
assign w3751 = w3748 & w3750;
assign w3752 = ~w3748 & ~w3750;
assign w3753 = ~w3751 & ~w3752;
assign w3754 = ~pi31 & pi33;
assign w3755 = ~w3530 & ~w3754;
assign w3756 = pi28 & w56;
assign w3757 = ~pi36 & pi37;
assign w3758 = ~w55 & ~w3757;
assign w3759 = pi35 & pi37;
assign w3760 = pi27 & ~w3759;
assign w3761 = ~w3758 & w3760;
assign w3762 = ~w3756 & ~w3761;
assign w3763 = pi37 & ~w3762;
assign w3764 = ~pi37 & w3762;
assign w3765 = ~w3763 & ~w3764;
assign w3766 = pi30 & w8;
assign w3767 = pi29 & ~w379;
assign w3768 = ~w378 & w3767;
assign w3769 = ~w3766 & ~w3768;
assign w3770 = pi35 & ~w3769;
assign w3771 = ~pi35 & w3769;
assign w3772 = ~w3770 & ~w3771;
assign w3773 = w3765 & w3772;
assign w3774 = ~w3765 & ~w3772;
assign w3775 = ~w3773 & ~w3774;
assign w3776 = w3755 & ~w3775;
assign w3777 = ~w3755 & w3775;
assign w3778 = ~w3776 & ~w3777;
assign w3779 = (~w3547 & ~w3549) | (~w3547 & w7628) | (~w3549 & w7628);
assign w3780 = ~w3778 & ~w3779;
assign w3781 = w3778 & w3779;
assign w3782 = ~w3780 & ~w3781;
assign w3783 = pi26 & w119;
assign w3784 = pi25 & ~w1634;
assign w3785 = ~w1633 & w3784;
assign w3786 = ~w3783 & ~w3785;
assign w3787 = pi39 & ~w3786;
assign w3788 = ~pi39 & w3786;
assign w3789 = ~w3787 & ~w3788;
assign w3790 = pi22 & w355;
assign w3791 = (pi43 & ~w353) | (pi43 & w8579) | (~w353 & w8579);
assign w3792 = pi21 & w354;
assign w3793 = ~w3790 & w8580;
assign w3794 = pi43 & w3790;
assign w3795 = ~w3793 & ~w3794;
assign w3796 = ~w3789 & ~w3795;
assign w3797 = w3789 & w3795;
assign w3798 = ~w3796 & ~w3797;
assign w3799 = pi24 & w217;
assign w3800 = (pi41 & ~w215) | (pi41 & w8581) | (~w215 & w8581);
assign w3801 = pi23 & w216;
assign w3802 = ~w3799 & w8582;
assign w3803 = pi41 & w3799;
assign w3804 = ~w3802 & ~w3803;
assign w3805 = w3798 & ~w3804;
assign w3806 = ~w3798 & w3804;
assign w3807 = ~w3805 & ~w3806;
assign w3808 = w3782 & ~w3807;
assign w3809 = ~w3782 & w3807;
assign w3810 = ~w3808 & ~w3809;
assign w3811 = w3753 & ~w3810;
assign w3812 = ~w3753 & w3810;
assign w3813 = ~w3811 & ~w3812;
assign w3814 = w3713 & ~w3813;
assign w3815 = ~w3713 & w3813;
assign w3816 = ~w3814 & ~w3815;
assign w3817 = w3662 & w3816;
assign w3818 = ~w3662 & ~w3816;
assign w3819 = ~w3817 & ~w3818;
assign w3820 = w3625 & ~w3819;
assign w3821 = ~w3625 & w3819;
assign w3822 = ~w3820 & ~w3821;
assign w3823 = ~w3620 & ~w3822;
assign w3824 = w3620 & w3822;
assign w3825 = ~w3823 & ~w3824;
assign w3826 = ~w3619 & w8583;
assign w3827 = (~w3825 & w3619) | (~w3825 & w8584) | (w3619 & w8584);
assign w3828 = ~w3826 & ~w3827;
assign w3829 = (~w3623 & ~w3625) | (~w3623 & w8585) | (~w3625 & w8585);
assign w3830 = ~w3651 & ~w3656;
assign w3831 = ~w3660 & ~w3816;
assign w3832 = (w3830 & w3831) | (w3830 & w7629) | (w3831 & w7629);
assign w3833 = ~w3831 & w7630;
assign w3834 = ~w3832 & ~w3833;
assign w3835 = (~w3642 & ~w3644) | (~w3642 & w8586) | (~w3644 & w8586);
assign w3836 = pi06 & ~w2588;
assign w3837 = pi07 & w2390;
assign w3838 = (pi59 & w3836) | (pi59 & w8587) | (w3836 & w8587);
assign w3839 = ~w3836 & w8588;
assign w3840 = ~w3838 & ~w3839;
assign w3841 = pi02 & ~w3404;
assign w3842 = pi03 & w3186;
assign w3843 = (pi63 & w3841) | (pi63 & w7631) | (w3841 & w7631);
assign w3844 = ~w3841 & w7632;
assign w3845 = ~w3843 & ~w3844;
assign w3846 = pi04 & ~w2981;
assign w3847 = pi05 & w2932;
assign w3848 = (pi61 & w3846) | (pi61 & w7633) | (w3846 & w7633);
assign w3849 = ~w3846 & w7634;
assign w3850 = ~w3848 & ~w3849;
assign w3851 = w3845 & w3850;
assign w3852 = ~w3845 & ~w3850;
assign w3853 = ~w3851 & ~w3852;
assign w3854 = w3840 & w3853;
assign w3855 = ~w3840 & ~w3853;
assign w3856 = ~w3854 & ~w3855;
assign w3857 = ~w3835 & w3856;
assign w3858 = w3835 & ~w3856;
assign w3859 = ~w3857 & ~w3858;
assign w3860 = w3649 & ~w3859;
assign w3861 = ~w3649 & w3859;
assign w3862 = ~w3860 & ~w3861;
assign w3863 = (~w3666 & ~w3667) | (~w3666 & w8589) | (~w3667 & w8589);
assign w3864 = ~w3862 & w3863;
assign w3865 = w3862 & ~w3863;
assign w3866 = ~w3864 & ~w3865;
assign w3867 = ~w3712 & w3813;
assign w3868 = ~w3711 & ~w3867;
assign w3869 = ~w3867 & w8590;
assign w3870 = (~w3866 & w3867) | (~w3866 & w8591) | (w3867 & w8591);
assign w3871 = ~w3869 & ~w3870;
assign w3872 = (~w3752 & w3810) | (~w3752 & w8592) | (w3810 & w8592);
assign w3873 = (~w3718 & ~w3745) | (~w3718 & w8593) | (~w3745 & w8593);
assign w3874 = (~w3675 & ~w3702) | (~w3675 & w8594) | (~w3702 & w8594);
assign w3875 = w3873 & w3874;
assign w3876 = ~w3873 & ~w3874;
assign w3877 = ~w3875 & ~w3876;
assign w3878 = pi08 & ~w2206;
assign w3879 = pi09 & w2032;
assign w3880 = (pi57 & w3878) | (pi57 & w8595) | (w3878 & w8595);
assign w3881 = ~w3878 & w8596;
assign w3882 = ~w3880 & ~w3881;
assign w3883 = (~w3699 & ~w3684) | (~w3699 & w8597) | (~w3684 & w8597);
assign w3884 = ~w3883 & w7635;
assign w3885 = (~w3882 & w3883) | (~w3882 & w7636) | (w3883 & w7636);
assign w3886 = ~w3884 & ~w3885;
assign w3887 = pi15 & w1132;
assign w3888 = pi14 & ~w2419;
assign w3889 = ~w2418 & w3888;
assign w3890 = ~w3887 & ~w3889;
assign w3891 = pi51 & ~w3890;
assign w3892 = ~pi51 & w3890;
assign w3893 = ~w3891 & ~w3892;
assign w3894 = pi13 & w1393;
assign w3895 = (pi53 & ~w1391) | (pi53 & w8598) | (~w1391 & w8598);
assign w3896 = pi12 & w1392;
assign w3897 = ~w3894 & w8599;
assign w3898 = pi53 & w3894;
assign w3899 = ~w3897 & ~w3898;
assign w3900 = ~w3893 & ~w3899;
assign w3901 = w3893 & w3899;
assign w3902 = ~w3900 & ~w3901;
assign w3903 = pi11 & w1695;
assign w3904 = (pi55 & ~w1693) | (pi55 & w8600) | (~w1693 & w8600);
assign w3905 = pi10 & w1694;
assign w3906 = ~w3903 & w8601;
assign w3907 = pi55 & w3903;
assign w3908 = ~w3906 & ~w3907;
assign w3909 = w3902 & ~w3908;
assign w3910 = ~w3902 & w3908;
assign w3911 = ~w3909 & ~w3910;
assign w3912 = w3886 & ~w3911;
assign w3913 = ~w3886 & w3911;
assign w3914 = ~w3912 & ~w3913;
assign w3915 = w3877 & w3914;
assign w3916 = ~w3877 & ~w3914;
assign w3917 = ~w3915 & ~w3916;
assign w3918 = w3872 & w3917;
assign w3919 = ~w3872 & ~w3917;
assign w3920 = ~w3918 & ~w3919;
assign w3921 = (~w3742 & ~w3727) | (~w3742 & w8602) | (~w3727 & w8602);
assign w3922 = ~w3734 & ~w3921;
assign w3923 = (~w3804 & ~w3789) | (~w3804 & w8603) | (~w3789 & w8603);
assign w3924 = ~w3796 & ~w3923;
assign w3925 = w3922 & w3924;
assign w3926 = ~w3922 & ~w3924;
assign w3927 = ~w3925 & ~w3926;
assign w3928 = pi21 & w523;
assign w3929 = pi20 & ~w1570;
assign w3930 = ~w1569 & w3929;
assign w3931 = ~w3928 & ~w3930;
assign w3932 = pi45 & ~w3931;
assign w3933 = ~pi45 & w3931;
assign w3934 = ~w3932 & ~w3933;
assign w3935 = pi19 & w700;
assign w3936 = (pi47 & ~w698) | (pi47 & w8604) | (~w698 & w8604);
assign w3937 = pi18 & w699;
assign w3938 = ~w3935 & w8605;
assign w3939 = pi47 & w3935;
assign w3940 = ~w3938 & ~w3939;
assign w3941 = ~w3934 & ~w3940;
assign w3942 = w3934 & w3940;
assign w3943 = ~w3941 & ~w3942;
assign w3944 = pi17 & w909;
assign w3945 = (pi49 & ~w907) | (pi49 & w8606) | (~w907 & w8606);
assign w3946 = pi16 & w908;
assign w3947 = ~w3944 & w8607;
assign w3948 = pi49 & w3944;
assign w3949 = ~w3947 & ~w3948;
assign w3950 = w3943 & ~w3949;
assign w3951 = ~w3943 & w3949;
assign w3952 = ~w3950 & ~w3951;
assign w3953 = w3927 & w3952;
assign w3954 = ~w3927 & ~w3952;
assign w3955 = ~w3953 & ~w3954;
assign w3956 = ~w3780 & w3807;
assign w3957 = ~w3781 & ~w3956;
assign w3958 = w3955 & ~w3957;
assign w3959 = ~w3955 & w3957;
assign w3960 = ~w3958 & ~w3959;
assign w3961 = pi30 & ~w25;
assign w3962 = pi31 & ~w7;
assign w3963 = ~w6 & w3962;
assign w3964 = (pi35 & w3961) | (pi35 & w7637) | (w3961 & w7637);
assign w3965 = ~w3961 & w7638;
assign w3966 = ~w3964 & ~w3965;
assign w3967 = pi28 & ~w2332;
assign w3968 = pi29 & w56;
assign w3969 = (pi37 & w3967) | (pi37 & w7639) | (w3967 & w7639);
assign w3970 = ~w3967 & w7640;
assign w3971 = ~w3969 & ~w3970;
assign w3972 = w3966 & w3971;
assign w3973 = ~w3966 & ~w3971;
assign w3974 = ~w3972 & ~w3973;
assign w3975 = (~w3774 & ~w3775) | (~w3774 & w7641) | (~w3775 & w7641);
assign w3976 = pi26 & ~w167;
assign w3977 = pi27 & w119;
assign w3978 = (pi39 & w3976) | (pi39 & w7642) | (w3976 & w7642);
assign w3979 = ~w3976 & w7643;
assign w3980 = ~w3978 & ~w3979;
assign w3981 = pi23 & w355;
assign w3982 = pi22 & ~w792;
assign w3983 = ~w791 & w3982;
assign w3984 = ~w3981 & ~w3983;
assign w3985 = pi43 & ~w3984;
assign w3986 = ~pi43 & w3984;
assign w3987 = ~w3985 & ~w3986;
assign w3988 = pi25 & w217;
assign w3989 = pi24 & ~w802;
assign w3990 = ~w801 & w3989;
assign w3991 = ~w3988 & ~w3990;
assign w3992 = pi41 & ~w3991;
assign w3993 = ~pi41 & w3991;
assign w3994 = ~w3992 & ~w3993;
assign w3995 = w3987 & w3994;
assign w3996 = ~w3987 & ~w3994;
assign w3997 = ~w3995 & ~w3996;
assign w3998 = w3980 & ~w3997;
assign w3999 = ~w3980 & w3997;
assign w4000 = ~w3998 & ~w3999;
assign w4001 = w3975 & ~w4000;
assign w4002 = ~w3975 & w4000;
assign w4003 = ~w4001 & ~w4002;
assign w4004 = w3974 & w4003;
assign w4005 = ~w3974 & ~w4003;
assign w4006 = ~w4004 & ~w4005;
assign w4007 = w3960 & ~w4006;
assign w4008 = ~w3960 & w4006;
assign w4009 = ~w4007 & ~w4008;
assign w4010 = w3920 & ~w4009;
assign w4011 = ~w3920 & w4009;
assign w4012 = ~w4010 & ~w4011;
assign w4013 = w3871 & w4012;
assign w4014 = ~w3871 & ~w4012;
assign w4015 = ~w4013 & ~w4014;
assign w4016 = w3834 & w4015;
assign w4017 = ~w3834 & ~w4015;
assign w4018 = ~w4016 & ~w4017;
assign w4019 = ~w3829 & w4018;
assign w4020 = w3829 & ~w4018;
assign w4021 = ~w4019 & ~w4020;
assign w4022 = ~w3596 & ~w3824;
assign w4023 = w4021 & w9083;
assign w4024 = (w3619 & w8608) | (w3619 & w8609) | (w8608 & w8609);
assign w4025 = ~w4023 & ~w4024;
assign w4026 = (~w3832 & ~w3834) | (~w3832 & w8610) | (~w3834 & w8610);
assign w4027 = ~w3861 & ~w3865;
assign w4028 = ~w3870 & ~w4012;
assign w4029 = (~w4027 & w4028) | (~w4027 & w7644) | (w4028 & w7644);
assign w4030 = ~w4028 & w7645;
assign w4031 = ~w4029 & ~w4030;
assign w4032 = ~w3919 & w4009;
assign w4033 = (~w3851 & ~w3853) | (~w3851 & w8611) | (~w3853 & w8611);
assign w4034 = pi07 & ~w2588;
assign w4035 = pi08 & w2390;
assign w4036 = (pi59 & w4034) | (pi59 & w8612) | (w4034 & w8612);
assign w4037 = ~w4034 & w8613;
assign w4038 = ~w4036 & ~w4037;
assign w4039 = pi03 & ~w3404;
assign w4040 = pi04 & w3186;
assign w4041 = (pi63 & w4039) | (pi63 & w7646) | (w4039 & w7646);
assign w4042 = ~w4039 & w7647;
assign w4043 = ~w4041 & ~w4042;
assign w4044 = pi05 & ~w2981;
assign w4045 = pi06 & w2932;
assign w4046 = (pi61 & w4044) | (pi61 & w7648) | (w4044 & w7648);
assign w4047 = ~w4044 & w7649;
assign w4048 = ~w4046 & ~w4047;
assign w4049 = w4043 & w4048;
assign w4050 = ~w4043 & ~w4048;
assign w4051 = ~w4049 & ~w4050;
assign w4052 = w4038 & w4051;
assign w4053 = ~w4038 & ~w4051;
assign w4054 = ~w4052 & ~w4053;
assign w4055 = ~w4033 & w4054;
assign w4056 = w4033 & ~w4054;
assign w4057 = ~w4055 & ~w4056;
assign w4058 = w3857 & w4057;
assign w4059 = ~w3857 & ~w4057;
assign w4060 = ~w4058 & ~w4059;
assign w4061 = ~w3875 & ~w3914;
assign w4062 = ~w3876 & ~w4061;
assign w4063 = w4060 & w4062;
assign w4064 = ~w4060 & ~w4062;
assign w4065 = ~w4063 & ~w4064;
assign w4066 = (w4065 & w4032) | (w4065 & w7650) | (w4032 & w7650);
assign w4067 = ~w3918 & ~w4065;
assign w4068 = ~w4032 & w4067;
assign w4069 = ~w4066 & ~w4068;
assign w4070 = pi09 & ~w2206;
assign w4071 = pi10 & w2032;
assign w4072 = (pi57 & w4070) | (pi57 & w8614) | (w4070 & w8614);
assign w4073 = ~w4070 & w8615;
assign w4074 = ~w4072 & ~w4073;
assign w4075 = (~w3908 & ~w3893) | (~w3908 & w8616) | (~w3893 & w8616);
assign w4076 = ~w4075 & w7651;
assign w4077 = (~w4074 & w4075) | (~w4074 & w7652) | (w4075 & w7652);
assign w4078 = ~w4076 & ~w4077;
assign w4079 = pi16 & w1132;
assign w4080 = pi15 & ~w2419;
assign w4081 = ~w2418 & w4080;
assign w4082 = ~w4079 & ~w4081;
assign w4083 = pi51 & ~w4082;
assign w4084 = ~pi51 & w4082;
assign w4085 = ~w4083 & ~w4084;
assign w4086 = pi12 & w1695;
assign w4087 = (pi55 & ~w1693) | (pi55 & w8617) | (~w1693 & w8617);
assign w4088 = pi11 & w1694;
assign w4089 = ~w4086 & w8618;
assign w4090 = pi55 & w4086;
assign w4091 = ~w4089 & ~w4090;
assign w4092 = ~w4085 & ~w4091;
assign w4093 = w4085 & w4091;
assign w4094 = ~w4092 & ~w4093;
assign w4095 = pi14 & w1393;
assign w4096 = (pi53 & ~w1391) | (pi53 & w8619) | (~w1391 & w8619);
assign w4097 = pi13 & w1392;
assign w4098 = ~w4095 & w8620;
assign w4099 = pi53 & w4095;
assign w4100 = ~w4098 & ~w4099;
assign w4101 = w4094 & ~w4100;
assign w4102 = ~w4094 & w4100;
assign w4103 = ~w4101 & ~w4102;
assign w4104 = ~w4078 & ~w4103;
assign w4105 = w4078 & w4103;
assign w4106 = ~w4104 & ~w4105;
assign w4107 = (~w3925 & w3952) | (~w3925 & w8621) | (w3952 & w8621);
assign w4108 = (~w3885 & ~w3911) | (~w3885 & w7653) | (~w3911 & w7653);
assign w4109 = w4107 & ~w4108;
assign w4110 = ~w4107 & w4108;
assign w4111 = ~w4109 & ~w4110;
assign w4112 = w4106 & w4111;
assign w4113 = ~w4106 & ~w4111;
assign w4114 = ~w4112 & ~w4113;
assign w4115 = ~w3959 & w4006;
assign w4116 = ~w3958 & ~w4115;
assign w4117 = w4114 & ~w4116;
assign w4118 = ~w4114 & w4116;
assign w4119 = ~w4117 & ~w4118;
assign w4120 = ~w3980 & ~w3995;
assign w4121 = ~w3996 & ~w4120;
assign w4122 = (~w3949 & ~w3934) | (~w3949 & w8622) | (~w3934 & w8622);
assign w4123 = ~w3941 & ~w4122;
assign w4124 = w4121 & w4123;
assign w4125 = ~w4121 & ~w4123;
assign w4126 = ~w4124 & ~w4125;
assign w4127 = pi22 & w523;
assign w4128 = pi21 & ~w1570;
assign w4129 = ~w1569 & w4128;
assign w4130 = ~w4127 & ~w4129;
assign w4131 = pi45 & ~w4130;
assign w4132 = ~pi45 & w4130;
assign w4133 = ~w4131 & ~w4132;
assign w4134 = pi20 & w700;
assign w4135 = (pi47 & ~w698) | (pi47 & w8623) | (~w698 & w8623);
assign w4136 = pi19 & w699;
assign w4137 = ~w4134 & w8624;
assign w4138 = pi47 & w4134;
assign w4139 = ~w4137 & ~w4138;
assign w4140 = ~w4133 & ~w4139;
assign w4141 = w4133 & w4139;
assign w4142 = ~w4140 & ~w4141;
assign w4143 = pi18 & w909;
assign w4144 = (pi49 & ~w907) | (pi49 & w8625) | (~w907 & w8625);
assign w4145 = pi17 & w908;
assign w4146 = ~w4143 & w8626;
assign w4147 = pi49 & w4143;
assign w4148 = ~w4146 & ~w4147;
assign w4149 = w4142 & ~w4148;
assign w4150 = ~w4142 & w4148;
assign w4151 = ~w4149 & ~w4150;
assign w4152 = w4126 & ~w4151;
assign w4153 = ~w4126 & w4151;
assign w4154 = ~w4152 & ~w4153;
assign w4155 = (~w3974 & ~w4000) | (~w3974 & w7654) | (~w4000 & w7654);
assign w4156 = ~w4001 & ~w4155;
assign w4157 = ~w4154 & w4156;
assign w4158 = w4154 & ~w4156;
assign w4159 = ~w4157 & ~w4158;
assign w4160 = pi30 & w56;
assign w4161 = pi29 & ~w3759;
assign w4162 = ~w3758 & w4161;
assign w4163 = ~w4160 & ~w4162;
assign w4164 = (pi35 & w7) | (pi35 & w7655) | (w7 & w7655);
assign w4165 = pi31 & ~pi35;
assign w4166 = ~w6 & w4165;
assign w4167 = pi37 & ~w4166;
assign w4168 = ~w4164 & w4167;
assign w4169 = w4163 & ~w4168;
assign w4170 = ~pi37 & ~w4166;
assign w4171 = ~w4164 & w4170;
assign w4172 = ~w4163 & ~w4171;
assign w4173 = ~w4169 & ~w4172;
assign w4174 = ~w4164 & ~w4166;
assign w4175 = ~pi37 & ~w4163;
assign w4176 = (~w4174 & ~w4163) | (~w4174 & w7656) | (~w4163 & w7656);
assign w4177 = ~w4175 & w4176;
assign w4178 = ~w4173 & ~w4177;
assign w4179 = w3973 & ~w4178;
assign w4180 = ~w3973 & w4178;
assign w4181 = ~w4179 & ~w4180;
assign w4182 = pi28 & w119;
assign w4183 = pi27 & ~w1634;
assign w4184 = ~w1633 & w4183;
assign w4185 = ~w4182 & ~w4184;
assign w4186 = pi39 & ~w4185;
assign w4187 = ~pi39 & w4185;
assign w4188 = ~w4186 & ~w4187;
assign w4189 = pi24 & w355;
assign w4190 = (pi43 & ~w353) | (pi43 & w8627) | (~w353 & w8627);
assign w4191 = pi23 & w354;
assign w4192 = ~w4189 & w8628;
assign w4193 = pi43 & w4189;
assign w4194 = ~w4192 & ~w4193;
assign w4195 = ~w4188 & ~w4194;
assign w4196 = w4188 & w4194;
assign w4197 = ~w4195 & ~w4196;
assign w4198 = pi26 & w217;
assign w4199 = (pi41 & ~w215) | (pi41 & w8629) | (~w215 & w8629);
assign w4200 = pi25 & w216;
assign w4201 = ~w4198 & w8630;
assign w4202 = pi41 & w4198;
assign w4203 = ~w4201 & ~w4202;
assign w4204 = w4197 & ~w4203;
assign w4205 = ~w4197 & w4203;
assign w4206 = ~w4204 & ~w4205;
assign w4207 = w4181 & ~w4206;
assign w4208 = ~w4181 & w4206;
assign w4209 = ~w4207 & ~w4208;
assign w4210 = w4159 & w4209;
assign w4211 = ~w4159 & ~w4209;
assign w4212 = ~w4210 & ~w4211;
assign w4213 = w4119 & ~w4212;
assign w4214 = ~w4119 & w4212;
assign w4215 = ~w4213 & ~w4214;
assign w4216 = w4069 & ~w4215;
assign w4217 = ~w4069 & w4215;
assign w4218 = ~w4216 & ~w4217;
assign w4219 = w4031 & w4218;
assign w4220 = ~w4031 & ~w4218;
assign w4221 = ~w4219 & ~w4220;
assign w4222 = ~w4026 & ~w4221;
assign w4223 = w4026 & w4221;
assign w4224 = ~w4222 & ~w4223;
assign w4225 = ~w2968 & w3606;
assign w4226 = w2371 & w2381;
assign w4227 = w2372 & w4226;
assign w4228 = w4225 & w8631;
assign w4229 = w2381 & w7657;
assign w4230 = ~w2572 & w2965;
assign w4231 = ~w4229 & w4230;
assign w4232 = w4225 & ~w4231;
assign w4233 = ~w3823 & ~w4020;
assign w4234 = ~w4019 & ~w4233;
assign w4235 = ~w3614 & w7891;
assign w4236 = ~w4232 & w4235;
assign w4237 = ~w4228 & w4236;
assign w4238 = ~w4019 & w4022;
assign w4239 = ~w4234 & ~w4238;
assign w4240 = (~w4239 & ~w4236) | (~w4239 & w8632) | (~w4236 & w8632);
assign w4241 = (w4236 & w8633) | (w4236 & w8634) | (w8633 & w8634);
assign w4242 = ~w4224 & w4240;
assign w4243 = ~w4241 & ~w4242;
assign w4244 = ~w4058 & ~w4063;
assign w4245 = ~w4244 & ~w4066;
assign w4246 = (w4245 & w4215) | (w4245 & w8635) | (w4215 & w8635);
assign w4247 = (w4244 & w4032) | (w4244 & w8950) | (w4032 & w8950);
assign w4248 = ~w4215 & w4247;
assign w4249 = (w4032 & w8636) | (w4032 & w8637) | (w8636 & w8637);
assign w4250 = (~w4249 & w4215) | (~w4249 & w8951) | (w4215 & w8951);
assign w4251 = ~w4246 & w4250;
assign w4252 = ~w4118 & ~w4212;
assign w4253 = (~w4049 & ~w4051) | (~w4049 & w8638) | (~w4051 & w8638);
assign w4254 = pi08 & ~w2588;
assign w4255 = pi09 & w2390;
assign w4256 = (pi59 & w4254) | (pi59 & w8639) | (w4254 & w8639);
assign w4257 = ~w4254 & w8640;
assign w4258 = ~w4256 & ~w4257;
assign w4259 = pi04 & ~w3404;
assign w4260 = pi05 & w3186;
assign w4261 = (pi63 & w4259) | (pi63 & w7658) | (w4259 & w7658);
assign w4262 = ~w4259 & w7659;
assign w4263 = ~w4261 & ~w4262;
assign w4264 = pi06 & ~w2981;
assign w4265 = pi07 & w2932;
assign w4266 = (pi61 & w4264) | (pi61 & w7660) | (w4264 & w7660);
assign w4267 = ~w4264 & w7661;
assign w4268 = ~w4266 & ~w4267;
assign w4269 = w4263 & w4268;
assign w4270 = ~w4263 & ~w4268;
assign w4271 = ~w4269 & ~w4270;
assign w4272 = w4258 & w4271;
assign w4273 = ~w4258 & ~w4271;
assign w4274 = ~w4272 & ~w4273;
assign w4275 = ~w4253 & w4274;
assign w4276 = w4253 & ~w4274;
assign w4277 = ~w4275 & ~w4276;
assign w4278 = w4055 & w4277;
assign w4279 = ~w4055 & ~w4277;
assign w4280 = ~w4278 & ~w4279;
assign w4281 = ~w4106 & ~w4109;
assign w4282 = ~w4110 & ~w4281;
assign w4283 = w4280 & ~w4282;
assign w4284 = ~w4280 & w4282;
assign w4285 = ~w4283 & ~w4284;
assign w4286 = ~w4117 & w4285;
assign w4287 = ~w4252 & w4286;
assign w4288 = (~w4285 & w4252) | (~w4285 & w7662) | (w4252 & w7662);
assign w4289 = ~w4287 & ~w4288;
assign w4290 = pi10 & ~w2206;
assign w4291 = pi11 & w2032;
assign w4292 = (pi57 & w4290) | (pi57 & w7893) | (w4290 & w7893);
assign w4293 = ~w4290 & w7894;
assign w4294 = ~w4292 & ~w4293;
assign w4295 = (~w4100 & ~w4085) | (~w4100 & w8641) | (~w4085 & w8641);
assign w4296 = ~w4295 & w7663;
assign w4297 = (~w4294 & w4295) | (~w4294 & w7664) | (w4295 & w7664);
assign w4298 = ~w4296 & ~w4297;
assign w4299 = pi16 & ~w1260;
assign w4300 = pi17 & w1132;
assign w4301 = (pi51 & w4299) | (pi51 & w8642) | (w4299 & w8642);
assign w4302 = ~w4299 & w8643;
assign w4303 = ~w4301 & ~w4302;
assign w4304 = pi15 & w1393;
assign w4305 = (pi53 & ~w1391) | (pi53 & w8644) | (~w1391 & w8644);
assign w4306 = pi14 & w1392;
assign w4307 = ~w4304 & w8645;
assign w4308 = pi53 & w4304;
assign w4309 = ~w4307 & ~w4308;
assign w4310 = pi13 & w1695;
assign w4311 = (pi55 & ~w1693) | (pi55 & w8646) | (~w1693 & w8646);
assign w4312 = pi12 & w1694;
assign w4313 = ~w4310 & w8647;
assign w4314 = pi55 & w4310;
assign w4315 = ~w4313 & ~w4314;
assign w4316 = ~w4309 & ~w4315;
assign w4317 = w4309 & w4315;
assign w4318 = ~w4316 & ~w4317;
assign w4319 = ~w4303 & w4318;
assign w4320 = w4303 & ~w4318;
assign w4321 = ~w4319 & ~w4320;
assign w4322 = w4298 & w4321;
assign w4323 = ~w4298 & ~w4321;
assign w4324 = ~w4322 & ~w4323;
assign w4325 = ~w4077 & ~w4105;
assign w4326 = ~w4324 & w4325;
assign w4327 = w4324 & ~w4325;
assign w4328 = ~w4326 & ~w4327;
assign w4329 = (~w4124 & ~w4126) | (~w4124 & w8648) | (~w4126 & w8648);
assign w4330 = ~w4328 & w4329;
assign w4331 = w4328 & ~w4329;
assign w4332 = ~w4330 & ~w4331;
assign w4333 = (~w4180 & w4206) | (~w4180 & w7665) | (w4206 & w7665);
assign w4334 = pi31 & ~w54;
assign w4335 = ~pi37 & ~w55;
assign w4336 = ~w4334 & w4335;
assign w4337 = pi30 & w54;
assign w4338 = w386 & w4334;
assign w4339 = w55 & w7666;
assign w4340 = ~w4336 & ~w4337;
assign w4341 = ~w4338 & ~w4339;
assign w4342 = w4340 & w4341;
assign w4343 = w4173 & ~w4342;
assign w4344 = ~w4173 & w4342;
assign w4345 = ~w4343 & ~w4344;
assign w4346 = pi28 & ~w167;
assign w4347 = pi29 & w119;
assign w4348 = (pi39 & w4346) | (pi39 & w7667) | (w4346 & w7667);
assign w4349 = ~w4346 & w7668;
assign w4350 = ~w4348 & ~w4349;
assign w4351 = pi27 & w217;
assign w4352 = pi26 & ~w802;
assign w4353 = ~w801 & w4352;
assign w4354 = ~w4351 & ~w4353;
assign w4355 = pi41 & ~w4354;
assign w4356 = ~pi41 & w4354;
assign w4357 = ~w4355 & ~w4356;
assign w4358 = pi25 & w355;
assign w4359 = pi24 & ~w792;
assign w4360 = ~w791 & w4359;
assign w4361 = ~w4358 & ~w4360;
assign w4362 = pi43 & ~w4361;
assign w4363 = ~pi43 & w4361;
assign w4364 = ~w4362 & ~w4363;
assign w4365 = ~w4357 & ~w4364;
assign w4366 = w4357 & w4364;
assign w4367 = ~w4365 & ~w4366;
assign w4368 = w4350 & ~w4367;
assign w4369 = ~w4350 & w4367;
assign w4370 = ~w4368 & ~w4369;
assign w4371 = w4345 & ~w4370;
assign w4372 = ~w4345 & w4370;
assign w4373 = ~w4371 & ~w4372;
assign w4374 = w4333 & ~w4373;
assign w4375 = ~w4333 & w4373;
assign w4376 = ~w4374 & ~w4375;
assign w4377 = (~w4148 & ~w4133) | (~w4148 & w8649) | (~w4133 & w8649);
assign w4378 = ~w4140 & ~w4377;
assign w4379 = (~w4203 & ~w4188) | (~w4203 & w8650) | (~w4188 & w8650);
assign w4380 = ~w4195 & ~w4379;
assign w4381 = ~w4378 & ~w4380;
assign w4382 = w4378 & w4380;
assign w4383 = ~w4381 & ~w4382;
assign w4384 = pi22 & ~w612;
assign w4385 = pi23 & w523;
assign w4386 = (pi45 & w4384) | (pi45 & w7669) | (w4384 & w7669);
assign w4387 = ~w4384 & w7670;
assign w4388 = ~w4386 & ~w4387;
assign w4389 = pi21 & w700;
assign w4390 = pi20 & ~w2099;
assign w4391 = ~w2098 & w4390;
assign w4392 = ~w4389 & ~w4391;
assign w4393 = pi47 & ~w4392;
assign w4394 = ~pi47 & w4392;
assign w4395 = ~w4393 & ~w4394;
assign w4396 = pi19 & w909;
assign w4397 = pi18 & ~w2273;
assign w4398 = ~w2272 & w4397;
assign w4399 = ~w4396 & ~w4398;
assign w4400 = pi49 & ~w4399;
assign w4401 = ~pi49 & w4399;
assign w4402 = ~w4400 & ~w4401;
assign w4403 = ~w4395 & ~w4402;
assign w4404 = w4395 & w4402;
assign w4405 = ~w4403 & ~w4404;
assign w4406 = w4388 & ~w4405;
assign w4407 = ~w4388 & w4405;
assign w4408 = ~w4406 & ~w4407;
assign w4409 = ~w4383 & w4408;
assign w4410 = w4383 & ~w4408;
assign w4411 = ~w4409 & ~w4410;
assign w4412 = ~w4376 & w4411;
assign w4413 = w4376 & ~w4411;
assign w4414 = ~w4412 & ~w4413;
assign w4415 = (~w4209 & ~w4154) | (~w4209 & w7671) | (~w4154 & w7671);
assign w4416 = ~w4157 & ~w4415;
assign w4417 = w4414 & ~w4416;
assign w4418 = ~w4414 & w4416;
assign w4419 = ~w4417 & ~w4418;
assign w4420 = w4332 & w4419;
assign w4421 = ~w4332 & ~w4419;
assign w4422 = ~w4420 & ~w4421;
assign w4423 = w4289 & ~w4422;
assign w4424 = ~w4289 & w4422;
assign w4425 = ~w4423 & ~w4424;
assign w4426 = ~w4251 & w4425;
assign w4427 = w4251 & ~w4425;
assign w4428 = ~w4426 & ~w4427;
assign w4429 = (~w4030 & w4218) | (~w4030 & w8651) | (w4218 & w8651);
assign w4430 = w4428 & ~w4429;
assign w4431 = ~w4428 & w4429;
assign w4432 = ~w4430 & ~w4431;
assign w4433 = ~w4222 & ~w4239;
assign w4434 = (~w4223 & w4239) | (~w4223 & w8652) | (w4239 & w8652);
assign w4435 = (~w4236 & w8653) | (~w4236 & w8654) | (w8653 & w8654);
assign w4436 = w4432 & w4435;
assign w4437 = ~w4432 & ~w4435;
assign w4438 = ~w4436 & ~w4437;
assign w4439 = ~w4248 & w8655;
assign w4440 = (~w4439 & w4251) | (~w4439 & w8656) | (w4251 & w8656);
assign w4441 = (~w4269 & ~w4271) | (~w4269 & w8657) | (~w4271 & w8657);
assign w4442 = pi09 & ~w2588;
assign w4443 = pi10 & w2390;
assign w4444 = (pi59 & w4442) | (pi59 & w8658) | (w4442 & w8658);
assign w4445 = ~w4442 & w8659;
assign w4446 = ~w4444 & ~w4445;
assign w4447 = pi05 & ~w3404;
assign w4448 = pi06 & w3186;
assign w4449 = (pi63 & w4447) | (pi63 & w8660) | (w4447 & w8660);
assign w4450 = ~w4447 & w8661;
assign w4451 = ~w4449 & ~w4450;
assign w4452 = pi07 & ~w2981;
assign w4453 = pi08 & w2932;
assign w4454 = (pi61 & w4452) | (pi61 & w8662) | (w4452 & w8662);
assign w4455 = ~w4452 & w8663;
assign w4456 = ~w4454 & ~w4455;
assign w4457 = w4451 & w4456;
assign w4458 = ~w4451 & ~w4456;
assign w4459 = ~w4457 & ~w4458;
assign w4460 = w4446 & w4459;
assign w4461 = ~w4446 & ~w4459;
assign w4462 = ~w4460 & ~w4461;
assign w4463 = ~w4441 & w4462;
assign w4464 = w4441 & ~w4462;
assign w4465 = ~w4463 & ~w4464;
assign w4466 = w4275 & w4465;
assign w4467 = ~w4275 & ~w4465;
assign w4468 = ~w4466 & ~w4467;
assign w4469 = (~w4326 & ~w4328) | (~w4326 & w8664) | (~w4328 & w8664);
assign w4470 = w4468 & ~w4469;
assign w4471 = ~w4468 & w4469;
assign w4472 = ~w4470 & ~w4471;
assign w4473 = (~w4382 & ~w4383) | (~w4382 & w7672) | (~w4383 & w7672);
assign w4474 = (~w4297 & ~w4298) | (~w4297 & w8665) | (~w4298 & w8665);
assign w4475 = w4473 & ~w4474;
assign w4476 = ~w4473 & w4474;
assign w4477 = ~w4475 & ~w4476;
assign w4478 = (~w4316 & ~w4318) | (~w4316 & w8666) | (~w4318 & w8666);
assign w4479 = pi11 & ~w2206;
assign w4480 = pi12 & w2032;
assign w4481 = (pi57 & w4479) | (pi57 & w8667) | (w4479 & w8667);
assign w4482 = ~w4479 & w8668;
assign w4483 = ~w4481 & ~w4482;
assign w4484 = pi18 & w1132;
assign w4485 = pi17 & ~w2419;
assign w4486 = ~w2418 & w4485;
assign w4487 = ~w4484 & ~w4486;
assign w4488 = pi51 & ~w4487;
assign w4489 = ~pi51 & w4487;
assign w4490 = ~w4488 & ~w4489;
assign w4491 = pi16 & w1393;
assign w4492 = (pi53 & ~w1391) | (pi53 & w8669) | (~w1391 & w8669);
assign w4493 = pi15 & w1392;
assign w4494 = ~w4491 & w8670;
assign w4495 = pi53 & w4491;
assign w4496 = ~w4494 & ~w4495;
assign w4497 = ~w4490 & ~w4496;
assign w4498 = w4490 & w4496;
assign w4499 = ~w4497 & ~w4498;
assign w4500 = pi14 & w1695;
assign w4501 = (pi55 & ~w1693) | (pi55 & w8671) | (~w1693 & w8671);
assign w4502 = pi13 & w1694;
assign w4503 = ~w4500 & w8672;
assign w4504 = pi55 & w4500;
assign w4505 = ~w4503 & ~w4504;
assign w4506 = w4499 & ~w4505;
assign w4507 = ~w4499 & w4505;
assign w4508 = ~w4506 & ~w4507;
assign w4509 = ~w4483 & w4508;
assign w4510 = w4483 & ~w4508;
assign w4511 = ~w4509 & ~w4510;
assign w4512 = w4478 & ~w4511;
assign w4513 = ~w4478 & w4511;
assign w4514 = ~w4512 & ~w4513;
assign w4515 = w4477 & w4514;
assign w4516 = ~w4477 & ~w4514;
assign w4517 = ~w4515 & ~w4516;
assign w4518 = ~w4350 & ~w4366;
assign w4519 = ~w4365 & ~w4518;
assign w4520 = ~w4388 & ~w4404;
assign w4521 = ~w4403 & ~w4520;
assign w4522 = w4519 & w4521;
assign w4523 = ~w4519 & ~w4521;
assign w4524 = ~w4522 & ~w4523;
assign w4525 = pi24 & w523;
assign w4526 = pi23 & ~w1570;
assign w4527 = ~w1569 & w4526;
assign w4528 = ~w4525 & ~w4527;
assign w4529 = pi45 & ~w4528;
assign w4530 = ~pi45 & w4528;
assign w4531 = ~w4529 & ~w4530;
assign w4532 = pi20 & w909;
assign w4533 = (pi49 & ~w907) | (pi49 & w8673) | (~w907 & w8673);
assign w4534 = pi19 & w908;
assign w4535 = ~w4532 & w8674;
assign w4536 = pi49 & w4532;
assign w4537 = ~w4535 & ~w4536;
assign w4538 = ~w4531 & ~w4537;
assign w4539 = w4531 & w4537;
assign w4540 = ~w4538 & ~w4539;
assign w4541 = pi22 & w700;
assign w4542 = (pi47 & ~w698) | (pi47 & w8675) | (~w698 & w8675);
assign w4543 = pi21 & w699;
assign w4544 = ~w4541 & w8676;
assign w4545 = pi47 & w4541;
assign w4546 = ~w4544 & ~w4545;
assign w4547 = w4540 & ~w4546;
assign w4548 = ~w4540 & w4546;
assign w4549 = ~w4547 & ~w4548;
assign w4550 = w4524 & ~w4549;
assign w4551 = ~w4524 & w4549;
assign w4552 = ~w4550 & ~w4551;
assign w4553 = w4367 & w7673;
assign w4554 = ~w4344 & w4350;
assign w4555 = ~w4367 & w4554;
assign w4556 = ~w4343 & ~w4555;
assign w4557 = ~w4553 & w4556;
assign w4558 = pi28 & w217;
assign w4559 = (pi41 & ~w215) | (pi41 & w8677) | (~w215 & w8677);
assign w4560 = pi27 & w216;
assign w4561 = ~w4558 & w8678;
assign w4562 = pi41 & w4558;
assign w4563 = ~w4561 & ~w4562;
assign w4564 = pi26 & w355;
assign w4565 = (pi43 & ~w353) | (pi43 & w8679) | (~w353 & w8679);
assign w4566 = pi25 & w354;
assign w4567 = ~w4564 & w8680;
assign w4568 = pi43 & w4564;
assign w4569 = ~w4567 & ~w4568;
assign w4570 = ~w4563 & ~w4569;
assign w4571 = w4563 & w4569;
assign w4572 = ~w4570 & ~w4571;
assign w4573 = (~pi37 & w54) | (~pi37 & w8681) | (w54 & w8681);
assign w4574 = ~w55 & w8682;
assign w4575 = ~w4573 & ~w4574;
assign w4576 = w4342 & ~w4575;
assign w4577 = ~w4342 & w4575;
assign w4578 = ~w4576 & ~w4577;
assign w4579 = pi30 & w119;
assign w4580 = (pi39 & ~w117) | (pi39 & w8683) | (~w117 & w8683);
assign w4581 = pi29 & w118;
assign w4582 = ~w4579 & w8684;
assign w4583 = pi39 & w4579;
assign w4584 = ~w4582 & ~w4583;
assign w4585 = w4578 & w4584;
assign w4586 = ~w4578 & ~w4584;
assign w4587 = ~w4585 & ~w4586;
assign w4588 = w4572 & w4587;
assign w4589 = ~w4572 & ~w4587;
assign w4590 = ~w4588 & ~w4589;
assign w4591 = w4557 & ~w4590;
assign w4592 = ~w4557 & w4590;
assign w4593 = ~w4591 & ~w4592;
assign w4594 = ~w4552 & w4593;
assign w4595 = w4552 & ~w4593;
assign w4596 = ~w4594 & ~w4595;
assign w4597 = ~w4374 & w4411;
assign w4598 = ~w4375 & ~w4597;
assign w4599 = ~w4596 & ~w4598;
assign w4600 = w4596 & w4598;
assign w4601 = ~w4599 & ~w4600;
assign w4602 = w4517 & ~w4601;
assign w4603 = ~w4517 & w4601;
assign w4604 = ~w4602 & ~w4603;
assign w4605 = ~w4332 & ~w4418;
assign w4606 = ~w4417 & ~w4605;
assign w4607 = ~w4604 & ~w4606;
assign w4608 = w4604 & w4606;
assign w4609 = ~w4607 & ~w4608;
assign w4610 = w4472 & w4609;
assign w4611 = ~w4472 & ~w4609;
assign w4612 = ~w4610 & ~w4611;
assign w4613 = ~w4288 & w4422;
assign w4614 = ~w4278 & ~w4283;
assign w4615 = w4422 & w7674;
assign w4616 = ~w4278 & w4287;
assign w4617 = ~w4287 & ~w4614;
assign w4618 = ~w4616 & ~w4617;
assign w4619 = ~w4613 & ~w4618;
assign w4620 = ~w4615 & ~w4619;
assign w4621 = w4612 & ~w4620;
assign w4622 = ~w4612 & w4620;
assign w4623 = ~w4621 & ~w4622;
assign w4624 = w4440 & w4623;
assign w4625 = ~w4440 & ~w4623;
assign w4626 = ~w4624 & ~w4625;
assign w4627 = ~w3597 & w4233;
assign w4628 = w4238 & w4627;
assign w4629 = ~w4223 & w4628;
assign w4630 = ~w3602 & w7895;
assign w4631 = ~w4430 & ~w4434;
assign w4632 = w4626 & w9084;
assign w4633 = (w4630 & w8685) | (w4630 & w8686) | (w8685 & w8686);
assign w4634 = ~w4632 & ~w4633;
assign w4635 = ~w4614 & ~w4619;
assign w4636 = ~w4621 & ~w4635;
assign w4637 = w4609 & w7675;
assign w4638 = w4467 & w4469;
assign w4639 = ~w4608 & w4638;
assign w4640 = (~w4466 & w4469) | (~w4466 & w8687) | (w4469 & w8687);
assign w4641 = w4607 & w4640;
assign w4642 = ~w4639 & ~w4641;
assign w4643 = w4608 & ~w4640;
assign w4644 = w4642 & ~w4643;
assign w4645 = (w4478 & ~w4508) | (w4478 & w8688) | (~w4508 & w8688);
assign w4646 = ~w4510 & ~w4645;
assign w4647 = pi12 & ~w2206;
assign w4648 = pi13 & w2032;
assign w4649 = (pi57 & w4647) | (pi57 & w8689) | (w4647 & w8689);
assign w4650 = ~w4647 & w8690;
assign w4651 = ~w4649 & ~w4650;
assign w4652 = (~w4505 & ~w4490) | (~w4505 & w8691) | (~w4490 & w8691);
assign w4653 = ~w4652 & w7676;
assign w4654 = (~w4651 & w4652) | (~w4651 & w7677) | (w4652 & w7677);
assign w4655 = ~w4653 & ~w4654;
assign w4656 = pi19 & w1132;
assign w4657 = pi18 & ~w1260;
assign w4658 = (pi51 & w4657) | (pi51 & w7678) | (w4657 & w7678);
assign w4659 = ~w4657 & w7679;
assign w4660 = ~w4658 & ~w4659;
assign w4661 = pi15 & w1695;
assign w4662 = (pi55 & ~w1693) | (pi55 & w8692) | (~w1693 & w8692);
assign w4663 = pi14 & w1694;
assign w4664 = ~w4661 & w8693;
assign w4665 = pi55 & w4661;
assign w4666 = ~w4664 & ~w4665;
assign w4667 = pi17 & w1393;
assign w4668 = (pi53 & ~w1391) | (pi53 & w8694) | (~w1391 & w8694);
assign w4669 = pi16 & w1392;
assign w4670 = ~w4667 & w8695;
assign w4671 = pi53 & w4667;
assign w4672 = ~w4670 & ~w4671;
assign w4673 = ~w4666 & ~w4672;
assign w4674 = w4666 & w4672;
assign w4675 = ~w4673 & ~w4674;
assign w4676 = w4660 & w4675;
assign w4677 = ~w4660 & ~w4675;
assign w4678 = ~w4676 & ~w4677;
assign w4679 = w4655 & w4678;
assign w4680 = ~w4655 & ~w4678;
assign w4681 = ~w4679 & ~w4680;
assign w4682 = w4646 & ~w4681;
assign w4683 = ~w4646 & w4681;
assign w4684 = ~w4682 & ~w4683;
assign w4685 = (~w4522 & ~w4524) | (~w4522 & w8696) | (~w4524 & w8696);
assign w4686 = w4684 & ~w4685;
assign w4687 = ~w4684 & w4685;
assign w4688 = ~w4686 & ~w4687;
assign w4689 = ~w4577 & ~w4584;
assign w4690 = ~w4572 & w4585;
assign w4691 = (~w4576 & ~w4572) | (~w4576 & w7680) | (~w4572 & w7680);
assign w4692 = ~w4690 & w4691;
assign w4693 = pi30 & ~w1634;
assign w4694 = ~w1633 & w4693;
assign w4695 = pi31 & ~w118;
assign w4696 = ~w117 & w4695;
assign w4697 = ~w4694 & ~w4696;
assign w4698 = pi39 & ~w4697;
assign w4699 = ~pi39 & w4697;
assign w4700 = ~w4698 & ~w4699;
assign w4701 = pi27 & w355;
assign w4702 = (pi43 & ~w353) | (pi43 & w8697) | (~w353 & w8697);
assign w4703 = pi26 & w354;
assign w4704 = ~w4701 & w8698;
assign w4705 = w355 & w9052;
assign w4706 = ~w4704 & ~w4705;
assign w4707 = ~w4700 & ~w4706;
assign w4708 = w4700 & w4706;
assign w4709 = ~w4707 & ~w4708;
assign w4710 = pi29 & w217;
assign w4711 = (pi41 & ~w215) | (pi41 & w8699) | (~w215 & w8699);
assign w4712 = pi28 & w216;
assign w4713 = ~w4710 & w8700;
assign w4714 = w217 & w9053;
assign w4715 = ~w4713 & ~w4714;
assign w4716 = w4709 & ~w4715;
assign w4717 = ~w4709 & w4715;
assign w4718 = ~w4716 & ~w4717;
assign w4719 = w4692 & ~w4718;
assign w4720 = ~w4692 & w4718;
assign w4721 = ~w4719 & ~w4720;
assign w4722 = ~w4571 & ~w4584;
assign w4723 = ~w4570 & ~w4722;
assign w4724 = (~w4546 & ~w4531) | (~w4546 & w8701) | (~w4531 & w8701);
assign w4725 = ~w4538 & ~w4724;
assign w4726 = ~w4723 & ~w4725;
assign w4727 = w4723 & w4725;
assign w4728 = ~w4726 & ~w4727;
assign w4729 = pi25 & w523;
assign w4730 = pi24 & ~w1570;
assign w4731 = ~w1569 & w4730;
assign w4732 = ~w4729 & ~w4731;
assign w4733 = pi45 & ~w4732;
assign w4734 = ~pi45 & w4732;
assign w4735 = ~w4733 & ~w4734;
assign w4736 = pi21 & w909;
assign w4737 = (pi49 & ~w907) | (pi49 & w8702) | (~w907 & w8702);
assign w4738 = pi20 & w908;
assign w4739 = ~w4736 & w8703;
assign w4740 = w909 & w9054;
assign w4741 = ~w4739 & ~w4740;
assign w4742 = ~w4735 & ~w4741;
assign w4743 = w4735 & w4741;
assign w4744 = ~w4742 & ~w4743;
assign w4745 = pi23 & w700;
assign w4746 = (pi47 & ~w698) | (pi47 & w8704) | (~w698 & w8704);
assign w4747 = pi22 & w699;
assign w4748 = ~w4745 & w8705;
assign w4749 = w700 & w9055;
assign w4750 = ~w4748 & ~w4749;
assign w4751 = w4744 & ~w4750;
assign w4752 = ~w4744 & w4750;
assign w4753 = ~w4751 & ~w4752;
assign w4754 = w4728 & ~w4753;
assign w4755 = ~w4728 & w4753;
assign w4756 = ~w4754 & ~w4755;
assign w4757 = w4721 & ~w4756;
assign w4758 = ~w4721 & w4756;
assign w4759 = ~w4757 & ~w4758;
assign w4760 = ~w4591 & ~w4594;
assign w4761 = w4759 & ~w4760;
assign w4762 = ~w4759 & w4760;
assign w4763 = ~w4761 & ~w4762;
assign w4764 = w4688 & w4763;
assign w4765 = ~w4688 & ~w4763;
assign w4766 = ~w4764 & ~w4765;
assign w4767 = (~w4457 & ~w4459) | (~w4457 & w8706) | (~w4459 & w8706);
assign w4768 = pi10 & ~w2588;
assign w4769 = pi11 & w2390;
assign w4770 = (pi59 & w4768) | (pi59 & w8707) | (w4768 & w8707);
assign w4771 = ~w4768 & w8708;
assign w4772 = ~w4770 & ~w4771;
assign w4773 = pi06 & ~w3404;
assign w4774 = pi07 & w3186;
assign w4775 = (pi63 & w4773) | (pi63 & w8709) | (w4773 & w8709);
assign w4776 = ~w4773 & w8710;
assign w4777 = ~w4775 & ~w4776;
assign w4778 = pi08 & ~w2981;
assign w4779 = pi09 & w2932;
assign w4780 = (pi61 & w4778) | (pi61 & w8711) | (w4778 & w8711);
assign w4781 = ~w4778 & w8712;
assign w4782 = ~w4780 & ~w4781;
assign w4783 = w4777 & w4782;
assign w4784 = ~w4777 & ~w4782;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = w4772 & w4785;
assign w4787 = ~w4772 & ~w4785;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = ~w4767 & w4788;
assign w4790 = w4767 & ~w4788;
assign w4791 = ~w4789 & ~w4790;
assign w4792 = w4463 & w4791;
assign w4793 = ~w4463 & ~w4791;
assign w4794 = ~w4792 & ~w4793;
assign w4795 = ~w4515 & w8713;
assign w4796 = (~w4794 & w4515) | (~w4794 & w8714) | (w4515 & w8714);
assign w4797 = ~w4795 & ~w4796;
assign w4798 = (~w4599 & ~w4601) | (~w4599 & w7681) | (~w4601 & w7681);
assign w4799 = w4797 & ~w4798;
assign w4800 = ~w4797 & w4798;
assign w4801 = ~w4799 & ~w4800;
assign w4802 = w4766 & ~w4801;
assign w4803 = ~w4766 & w4801;
assign w4804 = ~w4802 & ~w4803;
assign w4805 = (~w4804 & ~w4644) | (~w4804 & w7682) | (~w4644 & w7682);
assign w4806 = w4644 & w7683;
assign w4807 = ~w4805 & ~w4806;
assign w4808 = w4636 & w4807;
assign w4809 = ~w4636 & ~w4807;
assign w4810 = ~w4808 & ~w4809;
assign w4811 = w4432 & w4626;
assign w4812 = w4626 & w9056;
assign w4813 = w4628 & w4812;
assign w4814 = (w4813 & w3602) | (w4813 & w7684) | (w3602 & w7684);
assign w4815 = w4626 & w8952;
assign w4816 = ~w4628 & w4811;
assign w4817 = w4433 & w4816;
assign w4818 = ~w4431 & ~w4624;
assign w4819 = ~w4625 & ~w4818;
assign w4820 = ~w4817 & w7896;
assign w4821 = ~w4814 & w4820;
assign w4822 = (w4810 & w4814) | (w4810 & w8715) | (w4814 & w8715);
assign w4823 = ~w4814 & w8716;
assign w4824 = ~w4822 & ~w4823;
assign w4825 = w4640 & ~w4642;
assign w4826 = ~w4806 & ~w4825;
assign w4827 = ~w4792 & ~w4795;
assign w4828 = ~w4766 & ~w4799;
assign w4829 = ~w4828 & w7897;
assign w4830 = (w4827 & w4828) | (w4827 & w7898) | (w4828 & w7898);
assign w4831 = ~w4829 & ~w4830;
assign w4832 = (~w4762 & ~w4763) | (~w4762 & w8717) | (~w4763 & w8717);
assign w4833 = (~w4654 & w4678) | (~w4654 & w7685) | (w4678 & w7685);
assign w4834 = (~w4726 & ~w4753) | (~w4726 & w8718) | (~w4753 & w8718);
assign w4835 = ~w4833 & ~w4834;
assign w4836 = w4833 & w4834;
assign w4837 = ~w4835 & ~w4836;
assign w4838 = pi13 & ~w2206;
assign w4839 = pi14 & w2032;
assign w4840 = (pi57 & w4838) | (pi57 & w8719) | (w4838 & w8719);
assign w4841 = ~w4838 & w8720;
assign w4842 = ~w4840 & ~w4841;
assign w4843 = ~w4660 & ~w4674;
assign w4844 = ~w4843 & w7686;
assign w4845 = (~w4842 & w4843) | (~w4842 & w8721) | (w4843 & w8721);
assign w4846 = ~w4844 & ~w4845;
assign w4847 = pi20 & w1132;
assign w4848 = pi19 & ~w2419;
assign w4849 = ~w2418 & w4848;
assign w4850 = ~w4847 & ~w4849;
assign w4851 = pi51 & ~w4850;
assign w4852 = ~pi51 & w4850;
assign w4853 = ~w4851 & ~w4852;
assign w4854 = pi18 & w1393;
assign w4855 = (pi53 & ~w1391) | (pi53 & w8722) | (~w1391 & w8722);
assign w4856 = pi17 & w1392;
assign w4857 = ~w4854 & w8723;
assign w4858 = pi53 & w4854;
assign w4859 = ~w4857 & ~w4858;
assign w4860 = ~w4853 & ~w4859;
assign w4861 = w4853 & w4859;
assign w4862 = ~w4860 & ~w4861;
assign w4863 = pi16 & w1695;
assign w4864 = (pi55 & ~w1693) | (pi55 & w8724) | (~w1693 & w8724);
assign w4865 = pi15 & w1694;
assign w4866 = ~w4863 & w8725;
assign w4867 = pi55 & w4863;
assign w4868 = ~w4866 & ~w4867;
assign w4869 = w4862 & ~w4868;
assign w4870 = ~w4862 & w4868;
assign w4871 = ~w4869 & ~w4870;
assign w4872 = w4846 & ~w4871;
assign w4873 = ~w4846 & w4871;
assign w4874 = ~w4872 & ~w4873;
assign w4875 = ~w4837 & ~w4874;
assign w4876 = w4837 & w4874;
assign w4877 = ~w4875 & ~w4876;
assign w4878 = pi30 & w217;
assign w4879 = (pi41 & ~w215) | (pi41 & w8726) | (~w215 & w8726);
assign w4880 = pi29 & w216;
assign w4881 = ~w4878 & w8727;
assign w4882 = w217 & w9057;
assign w4883 = ~w4881 & ~w4882;
assign w4884 = pi28 & w355;
assign w4885 = (pi43 & ~w353) | (pi43 & w8728) | (~w353 & w8728);
assign w4886 = pi27 & w354;
assign w4887 = ~w4884 & w8729;
assign w4888 = w355 & w9058;
assign w4889 = ~w4887 & ~w4888;
assign w4890 = ~w4883 & ~w4889;
assign w4891 = w4883 & w4889;
assign w4892 = ~w4890 & ~w4891;
assign w4893 = (pi39 & w118) | (pi39 & w8730) | (w118 & w8730);
assign w4894 = pi31 & ~pi39;
assign w4895 = ~w117 & w4894;
assign w4896 = ~w4893 & ~w4895;
assign w4897 = ~w4892 & w4896;
assign w4898 = w4892 & ~w4896;
assign w4899 = ~w4897 & ~w4898;
assign w4900 = ~w4718 & ~w4899;
assign w4901 = w4718 & w4899;
assign w4902 = ~w4900 & ~w4901;
assign w4903 = (~w4750 & ~w4735) | (~w4750 & w8731) | (~w4735 & w8731);
assign w4904 = ~w4742 & ~w4903;
assign w4905 = (~w4715 & ~w4700) | (~w4715 & w8732) | (~w4700 & w8732);
assign w4906 = ~w4707 & ~w4905;
assign w4907 = w4904 & w4906;
assign w4908 = ~w4904 & ~w4906;
assign w4909 = ~w4907 & ~w4908;
assign w4910 = pi26 & w523;
assign w4911 = pi25 & ~w1570;
assign w4912 = ~w1569 & w4911;
assign w4913 = ~w4910 & ~w4912;
assign w4914 = pi45 & ~w4913;
assign w4915 = ~pi45 & w4913;
assign w4916 = ~w4914 & ~w4915;
assign w4917 = pi24 & w700;
assign w4918 = (pi47 & ~w698) | (pi47 & w8733) | (~w698 & w8733);
assign w4919 = pi23 & w699;
assign w4920 = ~w4917 & w8734;
assign w4921 = w700 & w9059;
assign w4922 = ~w4920 & ~w4921;
assign w4923 = ~w4916 & ~w4922;
assign w4924 = w4916 & w4922;
assign w4925 = ~w4923 & ~w4924;
assign w4926 = pi22 & w909;
assign w4927 = (pi49 & ~w907) | (pi49 & w8735) | (~w907 & w8735);
assign w4928 = pi21 & w908;
assign w4929 = ~w4926 & w8736;
assign w4930 = w909 & w9060;
assign w4931 = ~w4929 & ~w4930;
assign w4932 = w4925 & ~w4931;
assign w4933 = ~w4925 & w4931;
assign w4934 = ~w4932 & ~w4933;
assign w4935 = w4909 & ~w4934;
assign w4936 = ~w4909 & w4934;
assign w4937 = ~w4935 & ~w4936;
assign w4938 = w4902 & w4937;
assign w4939 = ~w4902 & ~w4937;
assign w4940 = ~w4938 & ~w4939;
assign w4941 = (~w4719 & w4756) | (~w4719 & w7687) | (w4756 & w7687);
assign w4942 = w4940 & w4941;
assign w4943 = ~w4940 & ~w4941;
assign w4944 = ~w4942 & ~w4943;
assign w4945 = w4877 & ~w4944;
assign w4946 = ~w4877 & w4944;
assign w4947 = ~w4945 & ~w4946;
assign w4948 = w4832 & w4947;
assign w4949 = ~w4832 & ~w4947;
assign w4950 = ~w4948 & ~w4949;
assign w4951 = (~w4683 & ~w4684) | (~w4683 & w8737) | (~w4684 & w8737);
assign w4952 = (~w4783 & ~w4785) | (~w4783 & w8738) | (~w4785 & w8738);
assign w4953 = pi11 & ~w2588;
assign w4954 = pi12 & w2390;
assign w4955 = (pi59 & w4953) | (pi59 & w8739) | (w4953 & w8739);
assign w4956 = ~w4953 & w8740;
assign w4957 = ~w4955 & ~w4956;
assign w4958 = pi07 & ~w3404;
assign w4959 = pi08 & w3186;
assign w4960 = (pi63 & w4958) | (pi63 & w8741) | (w4958 & w8741);
assign w4961 = ~w4958 & w8742;
assign w4962 = ~w4960 & ~w4961;
assign w4963 = pi09 & ~w2981;
assign w4964 = pi10 & w2932;
assign w4965 = (pi61 & w4963) | (pi61 & w8743) | (w4963 & w8743);
assign w4966 = ~w4963 & w8744;
assign w4967 = ~w4965 & ~w4966;
assign w4968 = w4962 & w4967;
assign w4969 = ~w4962 & ~w4967;
assign w4970 = ~w4968 & ~w4969;
assign w4971 = w4957 & w4970;
assign w4972 = ~w4957 & ~w4970;
assign w4973 = ~w4971 & ~w4972;
assign w4974 = ~w4952 & w4973;
assign w4975 = w4952 & ~w4973;
assign w4976 = ~w4974 & ~w4975;
assign w4977 = w4789 & w4976;
assign w4978 = ~w4789 & ~w4976;
assign w4979 = ~w4977 & ~w4978;
assign w4980 = ~w4951 & w4979;
assign w4981 = w4951 & ~w4979;
assign w4982 = ~w4980 & ~w4981;
assign w4983 = ~w4950 & w4982;
assign w4984 = w4950 & ~w4982;
assign w4985 = ~w4983 & ~w4984;
assign w4986 = w4831 & ~w4985;
assign w4987 = ~w4831 & w4985;
assign w4988 = ~w4986 & ~w4987;
assign w4989 = w4826 & w4988;
assign w4990 = ~w4826 & ~w4988;
assign w4991 = ~w4989 & ~w4990;
assign w4992 = (~w4809 & w4818) | (~w4809 & w7688) | (w4818 & w7688);
assign w4993 = (~w4808 & w4815) | (~w4808 & w7689) | (w4815 & w7689);
assign w4994 = (w7689 & w9061) | (w7689 & w9062) | (w9061 & w9062);
assign w4995 = w3598 & ~w4234;
assign w4996 = ~w3602 & w7690;
assign w4997 = w4811 & w7899;
assign w4998 = ~w4239 & w4997;
assign w4999 = w4997 & w8745;
assign w5000 = ~w4996 & w4999;
assign w5001 = (~w4994 & w4996) | (~w4994 & w7900) | (w4996 & w7900);
assign w5002 = ~w4991 & ~w4993;
assign w5003 = (w5002 & w4996) | (w5002 & w8746) | (w4996 & w8746);
assign w5004 = w5001 & ~w5003;
assign w5005 = (~w4829 & w4985) | (~w4829 & w7901) | (w4985 & w7901);
assign w5006 = ~w4949 & ~w4982;
assign w5007 = (~w4977 & w4951) | (~w4977 & w8747) | (w4951 & w8747);
assign w5008 = ~w4948 & ~w5007;
assign w5009 = ~w5006 & w5008;
assign w5010 = ~w4948 & w4982;
assign w5011 = ~w4949 & w5007;
assign w5012 = ~w5010 & w5011;
assign w5013 = ~w5009 & ~w5012;
assign w5014 = (~w4836 & ~w4837) | (~w4836 & w7691) | (~w4837 & w7691);
assign w5015 = (~w4968 & ~w4970) | (~w4968 & w8748) | (~w4970 & w8748);
assign w5016 = pi12 & ~w2588;
assign w5017 = pi13 & w2390;
assign w5018 = (pi59 & w5016) | (pi59 & w8749) | (w5016 & w8749);
assign w5019 = ~w5016 & w8750;
assign w5020 = ~w5018 & ~w5019;
assign w5021 = pi08 & ~w3404;
assign w5022 = pi09 & w3186;
assign w5023 = (pi63 & w5021) | (pi63 & w7902) | (w5021 & w7902);
assign w5024 = ~w5021 & w7903;
assign w5025 = ~w5023 & ~w5024;
assign w5026 = pi10 & ~w2981;
assign w5027 = pi11 & w2932;
assign w5028 = (pi61 & w5026) | (pi61 & w7904) | (w5026 & w7904);
assign w5029 = ~w5026 & w7905;
assign w5030 = ~w5028 & ~w5029;
assign w5031 = w5025 & w5030;
assign w5032 = ~w5025 & ~w5030;
assign w5033 = ~w5031 & ~w5032;
assign w5034 = w5020 & w5033;
assign w5035 = ~w5020 & ~w5033;
assign w5036 = ~w5034 & ~w5035;
assign w5037 = ~w5015 & w5036;
assign w5038 = w5015 & ~w5036;
assign w5039 = ~w5037 & ~w5038;
assign w5040 = w4974 & w5039;
assign w5041 = ~w4974 & ~w5039;
assign w5042 = ~w5040 & ~w5041;
assign w5043 = ~w5014 & w5042;
assign w5044 = w5014 & ~w5042;
assign w5045 = ~w5043 & ~w5044;
assign w5046 = w4877 & ~w4943;
assign w5047 = ~w4942 & ~w5046;
assign w5048 = w5045 & ~w5047;
assign w5049 = ~w5045 & w5047;
assign w5050 = ~w5048 & ~w5049;
assign w5051 = pi30 & ~w304;
assign w5052 = pi31 & ~w216;
assign w5053 = ~w215 & w5052;
assign w5054 = (pi41 & w5051) | (pi41 & w8751) | (w5051 & w8751);
assign w5055 = ~w5051 & w8752;
assign w5056 = ~w5054 & ~w5055;
assign w5057 = ~pi41 & w790;
assign w5058 = ~w439 & ~w5057;
assign w5059 = pi28 & ~w5058;
assign w5060 = pi29 & w355;
assign w5061 = (pi43 & w5059) | (pi43 & w8753) | (w5059 & w8753);
assign w5062 = ~w5059 & w8754;
assign w5063 = ~w5061 & ~w5062;
assign w5064 = w5056 & w5063;
assign w5065 = ~w5056 & ~w5063;
assign w5066 = ~w5064 & ~w5065;
assign w5067 = ~w4891 & ~w4896;
assign w5068 = ~w4890 & ~w5067;
assign w5069 = (~w4931 & ~w4916) | (~w4931 & w8755) | (~w4916 & w8755);
assign w5070 = ~w4923 & ~w5069;
assign w5071 = w5068 & w5070;
assign w5072 = ~w5068 & ~w5070;
assign w5073 = ~w5071 & ~w5072;
assign w5074 = pi27 & w523;
assign w5075 = pi26 & ~w1570;
assign w5076 = ~w1569 & w5075;
assign w5077 = ~w5074 & ~w5076;
assign w5078 = pi45 & ~w5077;
assign w5079 = ~pi45 & w5077;
assign w5080 = ~w5078 & ~w5079;
assign w5081 = pi25 & w700;
assign w5082 = (pi47 & ~w698) | (pi47 & w8756) | (~w698 & w8756);
assign w5083 = pi24 & w699;
assign w5084 = ~w5081 & w8757;
assign w5085 = w700 & w9063;
assign w5086 = ~w5084 & ~w5085;
assign w5087 = ~w5080 & ~w5086;
assign w5088 = w5080 & w5086;
assign w5089 = ~w5087 & ~w5088;
assign w5090 = pi23 & w909;
assign w5091 = (pi49 & ~w907) | (pi49 & w8758) | (~w907 & w8758);
assign w5092 = pi22 & w908;
assign w5093 = ~w5090 & w8759;
assign w5094 = w909 & w9064;
assign w5095 = ~w5093 & ~w5094;
assign w5096 = w5089 & ~w5095;
assign w5097 = ~w5089 & w5095;
assign w5098 = ~w5096 & ~w5097;
assign w5099 = w5073 & w5098;
assign w5100 = ~w5073 & ~w5098;
assign w5101 = ~w5099 & ~w5100;
assign w5102 = ~w5066 & ~w5101;
assign w5103 = w5066 & w5101;
assign w5104 = ~w5102 & ~w5103;
assign w5105 = (~w4900 & ~w4937) | (~w4900 & w7692) | (~w4937 & w7692);
assign w5106 = w5104 & ~w5105;
assign w5107 = ~w5104 & w5105;
assign w5108 = ~w5106 & ~w5107;
assign w5109 = (~w4845 & ~w4871) | (~w4845 & w8760) | (~w4871 & w8760);
assign w5110 = (~w4908 & ~w4934) | (~w4908 & w8761) | (~w4934 & w8761);
assign w5111 = w5109 & w5110;
assign w5112 = ~w5109 & ~w5110;
assign w5113 = ~w5111 & ~w5112;
assign w5114 = pi14 & ~w2206;
assign w5115 = pi15 & w2032;
assign w5116 = (pi57 & w5114) | (pi57 & w8762) | (w5114 & w8762);
assign w5117 = ~w5114 & w8763;
assign w5118 = ~w5116 & ~w5117;
assign w5119 = (~w4868 & ~w4853) | (~w4868 & w8764) | (~w4853 & w8764);
assign w5120 = ~w5119 & w7693;
assign w5121 = (~w5118 & w5119) | (~w5118 & w7906) | (w5119 & w7906);
assign w5122 = ~w5120 & ~w5121;
assign w5123 = pi21 & w1132;
assign w5124 = pi20 & ~w2419;
assign w5125 = ~w2418 & w5124;
assign w5126 = ~w5123 & ~w5125;
assign w5127 = pi51 & ~w5126;
assign w5128 = ~pi51 & w5126;
assign w5129 = ~w5127 & ~w5128;
assign w5130 = pi19 & w1393;
assign w5131 = (pi53 & ~w1391) | (pi53 & w8765) | (~w1391 & w8765);
assign w5132 = pi18 & w1392;
assign w5133 = ~w5130 & w8766;
assign w5134 = w1393 & w9065;
assign w5135 = ~w5133 & ~w5134;
assign w5136 = ~w5129 & ~w5135;
assign w5137 = w5129 & w5135;
assign w5138 = ~w5136 & ~w5137;
assign w5139 = pi17 & w1695;
assign w5140 = (pi55 & ~w1693) | (pi55 & w8767) | (~w1693 & w8767);
assign w5141 = pi16 & w1694;
assign w5142 = ~w5139 & w8768;
assign w5143 = w1695 & w9066;
assign w5144 = ~w5142 & ~w5143;
assign w5145 = w5138 & ~w5144;
assign w5146 = ~w5138 & w5144;
assign w5147 = ~w5145 & ~w5146;
assign w5148 = w5122 & ~w5147;
assign w5149 = ~w5122 & w5147;
assign w5150 = ~w5148 & ~w5149;
assign w5151 = ~w5113 & w5150;
assign w5152 = w5113 & ~w5150;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = w5108 & ~w5153;
assign w5155 = ~w5108 & w5153;
assign w5156 = ~w5154 & ~w5155;
assign w5157 = w5050 & w5156;
assign w5158 = ~w5050 & ~w5156;
assign w5159 = ~w5157 & ~w5158;
assign w5160 = w5013 & w5159;
assign w5161 = ~w5013 & ~w5159;
assign w5162 = ~w5160 & ~w5161;
assign w5163 = w5005 & ~w5162;
assign w5164 = ~w5005 & w5162;
assign w5165 = ~w5163 & ~w5164;
assign w5166 = w5165 & w9085;
assign w5167 = (w8025 & w8769) | (w8025 & w8770) | (w8769 & w8770);
assign w5168 = ~w5166 & ~w5167;
assign w5169 = (~w5009 & ~w5013) | (~w5009 & w7694) | (~w5013 & w7694);
assign w5170 = ~w5040 & ~w5043;
assign w5171 = ~w5048 & ~w5156;
assign w5172 = (w5170 & w5171) | (w5170 & w7695) | (w5171 & w7695);
assign w5173 = ~w5171 & w7696;
assign w5174 = ~w5172 & ~w5173;
assign w5175 = (~w5031 & ~w5033) | (~w5031 & w8771) | (~w5033 & w8771);
assign w5176 = pi13 & ~w2588;
assign w5177 = pi14 & w2390;
assign w5178 = (pi59 & w5176) | (pi59 & w8772) | (w5176 & w8772);
assign w5179 = ~w5176 & w8773;
assign w5180 = ~w5178 & ~w5179;
assign w5181 = pi09 & ~w3404;
assign w5182 = pi10 & w3186;
assign w5183 = (pi63 & w5181) | (pi63 & w7907) | (w5181 & w7907);
assign w5184 = ~w5181 & w7908;
assign w5185 = ~w5183 & ~w5184;
assign w5186 = pi11 & ~w2981;
assign w5187 = pi12 & w2932;
assign w5188 = (pi61 & w5186) | (pi61 & w7909) | (w5186 & w7909);
assign w5189 = ~w5186 & w7910;
assign w5190 = ~w5188 & ~w5189;
assign w5191 = w5185 & w5190;
assign w5192 = ~w5185 & ~w5190;
assign w5193 = ~w5191 & ~w5192;
assign w5194 = w5180 & w5193;
assign w5195 = ~w5180 & ~w5193;
assign w5196 = ~w5194 & ~w5195;
assign w5197 = ~w5175 & w5196;
assign w5198 = w5175 & ~w5196;
assign w5199 = ~w5197 & ~w5198;
assign w5200 = w5037 & w5199;
assign w5201 = ~w5037 & ~w5199;
assign w5202 = ~w5200 & ~w5201;
assign w5203 = (~w5112 & ~w5113) | (~w5112 & w7697) | (~w5113 & w7697);
assign w5204 = w5202 & w5203;
assign w5205 = ~w5202 & ~w5203;
assign w5206 = ~w5204 & ~w5205;
assign w5207 = (~w5106 & ~w5108) | (~w5106 & w7698) | (~w5108 & w7698);
assign w5208 = w5206 & ~w5207;
assign w5209 = ~w5206 & w5207;
assign w5210 = ~w5208 & ~w5209;
assign w5211 = (~w5121 & ~w5147) | (~w5121 & w7911) | (~w5147 & w7911);
assign w5212 = (~w5071 & w5098) | (~w5071 & w8774) | (w5098 & w8774);
assign w5213 = w5211 & ~w5212;
assign w5214 = ~w5211 & w5212;
assign w5215 = ~w5213 & ~w5214;
assign w5216 = pi15 & ~w2206;
assign w5217 = pi16 & w2032;
assign w5218 = (pi57 & w5216) | (pi57 & w8775) | (w5216 & w8775);
assign w5219 = ~w5216 & w8776;
assign w5220 = ~w5218 & ~w5219;
assign w5221 = (~w5144 & ~w5129) | (~w5144 & w8777) | (~w5129 & w8777);
assign w5222 = ~w5136 & ~w5221;
assign w5223 = ~w5221 & w7699;
assign w5224 = ~w5220 & ~w5222;
assign w5225 = ~w5223 & ~w5224;
assign w5226 = pi22 & w1132;
assign w5227 = pi21 & ~w2419;
assign w5228 = ~w2418 & w5227;
assign w5229 = ~w5226 & ~w5228;
assign w5230 = pi51 & ~w5229;
assign w5231 = ~pi51 & w5229;
assign w5232 = ~w5230 & ~w5231;
assign w5233 = pi20 & w1393;
assign w5234 = (pi53 & ~w1391) | (pi53 & w8778) | (~w1391 & w8778);
assign w5235 = pi19 & w1392;
assign w5236 = ~w5233 & w8779;
assign w5237 = w1393 & w9067;
assign w5238 = ~w5236 & ~w5237;
assign w5239 = ~w5232 & ~w5238;
assign w5240 = w5232 & w5238;
assign w5241 = ~w5239 & ~w5240;
assign w5242 = pi18 & w1695;
assign w5243 = (pi55 & ~w1693) | (pi55 & w8780) | (~w1693 & w8780);
assign w5244 = pi17 & w1694;
assign w5245 = ~w5242 & w8781;
assign w5246 = w1695 & w9068;
assign w5247 = ~w5245 & ~w5246;
assign w5248 = w5241 & ~w5247;
assign w5249 = ~w5241 & w5247;
assign w5250 = ~w5248 & ~w5249;
assign w5251 = w5225 & ~w5250;
assign w5252 = ~w5225 & w5250;
assign w5253 = ~w5251 & ~w5252;
assign w5254 = w5215 & ~w5253;
assign w5255 = ~w5215 & w5253;
assign w5256 = ~w5254 & ~w5255;
assign w5257 = (~w5095 & ~w5080) | (~w5095 & w8782) | (~w5080 & w8782);
assign w5258 = ~w5087 & ~w5257;
assign w5259 = w5065 & ~w5258;
assign w5260 = ~w5065 & w5258;
assign w5261 = ~w5259 & ~w5260;
assign w5262 = pi29 & ~w5058;
assign w5263 = pi30 & w355;
assign w5264 = (pi43 & w5262) | (pi43 & w8783) | (w5262 & w8783);
assign w5265 = ~w5262 & w8784;
assign w5266 = ~w5264 & ~w5265;
assign w5267 = (pi41 & w216) | (pi41 & w8785) | (w216 & w8785);
assign w5268 = pi31 & ~pi41;
assign w5269 = ~w215 & w5268;
assign w5270 = ~w5267 & ~w5269;
assign w5271 = ~w5266 & ~w5270;
assign w5272 = w5266 & w5270;
assign w5273 = ~w5271 & ~w5272;
assign w5274 = pi28 & w523;
assign w5275 = pi27 & ~w1570;
assign w5276 = ~w1569 & w5275;
assign w5277 = ~w5274 & ~w5276;
assign w5278 = pi45 & ~w5277;
assign w5279 = ~pi45 & w5277;
assign w5280 = ~w5278 & ~w5279;
assign w5281 = pi24 & w909;
assign w5282 = (pi49 & ~w907) | (pi49 & w8786) | (~w907 & w8786);
assign w5283 = pi23 & w908;
assign w5284 = ~w5281 & w8787;
assign w5285 = w909 & w9069;
assign w5286 = ~w5284 & ~w5285;
assign w5287 = ~w5280 & ~w5286;
assign w5288 = w5280 & w5286;
assign w5289 = ~w5287 & ~w5288;
assign w5290 = pi26 & w700;
assign w5291 = (pi47 & ~w698) | (pi47 & w8788) | (~w698 & w8788);
assign w5292 = pi25 & w699;
assign w5293 = ~w5290 & w8789;
assign w5294 = w700 & w9070;
assign w5295 = ~w5293 & ~w5294;
assign w5296 = w5289 & ~w5295;
assign w5297 = ~w5289 & w5295;
assign w5298 = ~w5296 & ~w5297;
assign w5299 = w5273 & ~w5298;
assign w5300 = ~w5273 & w5298;
assign w5301 = ~w5299 & ~w5300;
assign w5302 = w5261 & w5301;
assign w5303 = ~w5261 & ~w5301;
assign w5304 = ~w5302 & ~w5303;
assign w5305 = w5102 & w5304;
assign w5306 = ~w5102 & ~w5304;
assign w5307 = ~w5305 & ~w5306;
assign w5308 = ~w5256 & w5307;
assign w5309 = w5256 & ~w5307;
assign w5310 = ~w5308 & ~w5309;
assign w5311 = w5210 & w5310;
assign w5312 = ~w5210 & ~w5310;
assign w5313 = ~w5311 & ~w5312;
assign w5314 = ~w5174 & w5313;
assign w5315 = w5174 & ~w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = ~w5169 & ~w5316;
assign w5318 = w5169 & w5316;
assign w5319 = ~w5317 & ~w5318;
assign w5320 = w4991 & w5165;
assign w5321 = w4810 & w5320;
assign w5322 = w5320 & w7912;
assign w5323 = w4811 & w7913;
assign w5324 = w5322 & w5323;
assign w5325 = ~w3617 & w7914;
assign w5326 = w4811 & w7915;
assign w5327 = w5322 & w5326;
assign w5328 = (~w5327 & ~w3613) | (~w5327 & w7700) | (~w3613 & w7700);
assign w5329 = ~w5325 & w5328;
assign w5330 = ~w4989 & ~w5164;
assign w5331 = (~w5163 & w4989) | (~w5163 & w8790) | (w4989 & w8790);
assign w5332 = (~w4989 & ~w4812) | (~w4989 & w7701) | (~w4812 & w7701);
assign w5333 = ~w4993 & w5332;
assign w5334 = (w5320 & w4993) | (w5320 & w9071) | (w4993 & w9071);
assign w5335 = (~w5331 & w5333) | (~w5331 & w8791) | (w5333 & w8791);
assign w5336 = (w5319 & ~w5329) | (w5319 & w7916) | (~w5329 & w7916);
assign w5337 = w5329 & w8026;
assign w5338 = ~w5336 & ~w5337;
assign w5339 = (~w5305 & ~w5307) | (~w5305 & w8792) | (~w5307 & w8792);
assign w5340 = (~w5260 & w5298) | (~w5260 & w8793) | (w5298 & w8793);
assign w5341 = (~w5224 & ~w5250) | (~w5224 & w8794) | (~w5250 & w8794);
assign w5342 = ~w5340 & w5341;
assign w5343 = w5340 & ~w5341;
assign w5344 = ~w5342 & ~w5343;
assign w5345 = pi16 & ~w2206;
assign w5346 = pi17 & w2032;
assign w5347 = (pi57 & w5345) | (pi57 & w8795) | (w5345 & w8795);
assign w5348 = ~w5345 & w8796;
assign w5349 = ~w5347 & ~w5348;
assign w5350 = (~w5247 & ~w5232) | (~w5247 & w8797) | (~w5232 & w8797);
assign w5351 = ~w5239 & ~w5350;
assign w5352 = ~w5350 & w7702;
assign w5353 = ~w5349 & ~w5351;
assign w5354 = ~w5352 & ~w5353;
assign w5355 = pi23 & w1132;
assign w5356 = pi22 & ~w2419;
assign w5357 = ~w2418 & w5356;
assign w5358 = ~w5355 & ~w5357;
assign w5359 = pi51 & ~w5358;
assign w5360 = ~pi51 & w5358;
assign w5361 = ~w5359 & ~w5360;
assign w5362 = pi21 & w1393;
assign w5363 = (pi53 & ~w1391) | (pi53 & w8798) | (~w1391 & w8798);
assign w5364 = pi20 & w1392;
assign w5365 = ~w5362 & w8799;
assign w5366 = pi53 & w5362;
assign w5367 = ~w5365 & ~w5366;
assign w5368 = ~w5361 & ~w5367;
assign w5369 = w5361 & w5367;
assign w5370 = ~w5368 & ~w5369;
assign w5371 = pi19 & w1695;
assign w5372 = (pi55 & ~w1693) | (pi55 & w8800) | (~w1693 & w8800);
assign w5373 = pi18 & w1694;
assign w5374 = ~w5371 & w8801;
assign w5375 = pi55 & w5371;
assign w5376 = ~w5374 & ~w5375;
assign w5377 = w5370 & ~w5376;
assign w5378 = ~w5370 & w5376;
assign w5379 = ~w5377 & ~w5378;
assign w5380 = w5354 & ~w5379;
assign w5381 = ~w5354 & w5379;
assign w5382 = ~w5380 & ~w5381;
assign w5383 = w5344 & ~w5382;
assign w5384 = ~w5344 & w5382;
assign w5385 = ~w5383 & ~w5384;
assign w5386 = ~w5298 & w5261;
assign w5387 = (w5273 & w5261) | (w5273 & w5299) | (w5261 & w5299);
assign w5388 = ~w5386 & w5387;
assign w5389 = (~w5295 & ~w5280) | (~w5295 & w8802) | (~w5280 & w8802);
assign w5390 = ~w5287 & ~w5389;
assign w5391 = w5272 & w5390;
assign w5392 = ~w5272 & ~w5390;
assign w5393 = ~w5391 & ~w5392;
assign w5394 = pi28 & ~w612;
assign w5395 = pi29 & w523;
assign w5396 = (pi45 & w5394) | (pi45 & w8803) | (w5394 & w8803);
assign w5397 = ~w5394 & w8804;
assign w5398 = ~w5396 & ~w5397;
assign w5399 = pi25 & w909;
assign w5400 = (pi49 & ~w907) | (pi49 & w8805) | (~w907 & w8805);
assign w5401 = pi24 & w908;
assign w5402 = ~w5399 & w8806;
assign w5403 = w909 & w9072;
assign w5404 = ~w5402 & ~w5403;
assign w5405 = pi27 & w700;
assign w5406 = (pi47 & ~w698) | (pi47 & w8807) | (~w698 & w8807);
assign w5407 = pi26 & w699;
assign w5408 = ~w5405 & w8808;
assign w5409 = w700 & w9073;
assign w5410 = ~w5408 & ~w5409;
assign w5411 = w5404 & w5410;
assign w5412 = ~w5404 & ~w5410;
assign w5413 = ~w5411 & ~w5412;
assign w5414 = w5398 & w5413;
assign w5415 = ~w5398 & ~w5413;
assign w5416 = ~w5414 & ~w5415;
assign w5417 = pi30 & ~w5058;
assign w5418 = ~w438 & ~w790;
assign w5419 = pi31 & ~w5418;
assign w5420 = ~w5417 & ~w5419;
assign w5421 = (~w355 & w5058) | (~w355 & w8809) | (w5058 & w8809);
assign w5422 = pi31 & ~w5421;
assign w5423 = ~w5420 & ~w5422;
assign w5424 = pi31 & w355;
assign w5425 = ~w5419 & ~w5424;
assign w5426 = pi43 & ~w5425;
assign w5427 = ~pi43 & w5425;
assign w5428 = ~w5426 & ~w5427;
assign w5429 = ~w5423 & ~w5428;
assign w5430 = w5423 & w5428;
assign w5431 = ~w5429 & ~w5430;
assign w5432 = w5416 & ~w5431;
assign w5433 = ~w5416 & w5431;
assign w5434 = ~w5432 & ~w5433;
assign w5435 = w5393 & ~w5434;
assign w5436 = ~w5393 & w5434;
assign w5437 = ~w5435 & ~w5436;
assign w5438 = w5388 & ~w5437;
assign w5439 = ~w5388 & w5437;
assign w5440 = ~w5438 & ~w5439;
assign w5441 = ~w5385 & w5440;
assign w5442 = w5385 & ~w5440;
assign w5443 = ~w5441 & ~w5442;
assign w5444 = ~w5339 & w5443;
assign w5445 = w5339 & ~w5443;
assign w5446 = ~w5444 & ~w5445;
assign w5447 = (~w5191 & ~w5193) | (~w5191 & w8810) | (~w5193 & w8810);
assign w5448 = pi14 & ~w2588;
assign w5449 = pi15 & w2390;
assign w5450 = (pi59 & w5448) | (pi59 & w8811) | (w5448 & w8811);
assign w5451 = ~w5448 & w8812;
assign w5452 = ~w5450 & ~w5451;
assign w5453 = pi10 & ~w3404;
assign w5454 = pi11 & w3186;
assign w5455 = (pi63 & w5453) | (pi63 & w8813) | (w5453 & w8813);
assign w5456 = ~w5453 & w8814;
assign w5457 = ~w5455 & ~w5456;
assign w5458 = pi12 & ~w2981;
assign w5459 = pi13 & w2932;
assign w5460 = (pi61 & w5458) | (pi61 & w8815) | (w5458 & w8815);
assign w5461 = ~w5458 & w8816;
assign w5462 = ~w5460 & ~w5461;
assign w5463 = w5457 & w5462;
assign w5464 = ~w5457 & ~w5462;
assign w5465 = ~w5463 & ~w5464;
assign w5466 = w5452 & w5465;
assign w5467 = ~w5452 & ~w5465;
assign w5468 = ~w5466 & ~w5467;
assign w5469 = ~w5447 & w5468;
assign w5470 = w5447 & ~w5468;
assign w5471 = ~w5469 & ~w5470;
assign w5472 = w5197 & w5471;
assign w5473 = ~w5197 & ~w5471;
assign w5474 = ~w5472 & ~w5473;
assign w5475 = (~w5214 & ~w5215) | (~w5214 & w8817) | (~w5215 & w8817);
assign w5476 = w5474 & w5475;
assign w5477 = ~w5474 & ~w5475;
assign w5478 = ~w5476 & ~w5477;
assign w5479 = ~w5446 & ~w5478;
assign w5480 = w5446 & w5478;
assign w5481 = ~w5479 & ~w5480;
assign w5482 = ~w5207 & ~w5310;
assign w5483 = ~w5209 & ~w5482;
assign w5484 = ~w5310 & w7703;
assign w5485 = (~w5200 & ~w5203) | (~w5200 & w7917) | (~w5203 & w7917);
assign w5486 = (~w5485 & w5310) | (~w5485 & w7704) | (w5310 & w7704);
assign w5487 = ~w5484 & ~w5486;
assign w5488 = w5483 & ~w5487;
assign w5489 = ~w5483 & w5487;
assign w5490 = ~w5488 & ~w5489;
assign w5491 = w5481 & ~w5490;
assign w5492 = ~w5481 & w5490;
assign w5493 = ~w5491 & ~w5492;
assign w5494 = ~w5172 & ~w5315;
assign w5495 = w5493 & ~w5494;
assign w5496 = ~w5493 & w5494;
assign w5497 = ~w5495 & ~w5496;
assign w5498 = w5497 & w5336;
assign w5499 = w5317 & ~w5497;
assign w5500 = ~w5317 & w5497;
assign w5501 = ~w5499 & ~w5500;
assign w5502 = (w5329 & w8027) | (w5329 & w8028) | (w8027 & w8028);
assign w5503 = ~w5498 & ~w5502;
assign w5504 = w5485 & ~w5490;
assign w5505 = ~w5492 & ~w5504;
assign w5506 = w5446 & w7705;
assign w5507 = w5473 & ~w5475;
assign w5508 = ~w5444 & w5507;
assign w5509 = ~w5472 & ~w5476;
assign w5510 = w5445 & w5509;
assign w5511 = ~w5508 & ~w5510;
assign w5512 = w5444 & ~w5509;
assign w5513 = w5511 & ~w5512;
assign w5514 = ~w5506 & w5513;
assign w5515 = (~w5343 & ~w5344) | (~w5343 & w7706) | (~w5344 & w7706);
assign w5516 = (~w5463 & ~w5465) | (~w5463 & w8818) | (~w5465 & w8818);
assign w5517 = pi15 & ~w2588;
assign w5518 = pi16 & w2390;
assign w5519 = (pi59 & w5517) | (pi59 & w8819) | (w5517 & w8819);
assign w5520 = ~w5517 & w8820;
assign w5521 = ~w5519 & ~w5520;
assign w5522 = pi11 & ~w3404;
assign w5523 = pi12 & w3186;
assign w5524 = (pi63 & w5522) | (pi63 & w8821) | (w5522 & w8821);
assign w5525 = ~w5522 & w8822;
assign w5526 = ~w5524 & ~w5525;
assign w5527 = pi13 & ~w2981;
assign w5528 = pi14 & w2932;
assign w5529 = (pi61 & w5527) | (pi61 & w8823) | (w5527 & w8823);
assign w5530 = ~w5527 & w8824;
assign w5531 = ~w5529 & ~w5530;
assign w5532 = w5526 & w5531;
assign w5533 = ~w5526 & ~w5531;
assign w5534 = ~w5532 & ~w5533;
assign w5535 = w5521 & w5534;
assign w5536 = ~w5521 & ~w5534;
assign w5537 = ~w5535 & ~w5536;
assign w5538 = ~w5516 & w5537;
assign w5539 = w5516 & ~w5537;
assign w5540 = ~w5538 & ~w5539;
assign w5541 = w5469 & w5540;
assign w5542 = ~w5469 & ~w5540;
assign w5543 = ~w5541 & ~w5542;
assign w5544 = w5515 & w5543;
assign w5545 = ~w5515 & ~w5543;
assign w5546 = ~w5544 & ~w5545;
assign w5547 = ~w5438 & ~w5441;
assign w5548 = w5546 & ~w5547;
assign w5549 = ~w5546 & w5547;
assign w5550 = ~w5548 & ~w5549;
assign w5551 = (~w5353 & ~w5379) | (~w5353 & w8825) | (~w5379 & w8825);
assign w5552 = ~w5392 & w5416;
assign w5553 = ~w5391 & ~w5552;
assign w5554 = w5551 & ~w5553;
assign w5555 = ~w5551 & w5553;
assign w5556 = ~w5554 & ~w5555;
assign w5557 = pi17 & ~w2206;
assign w5558 = pi18 & w2032;
assign w5559 = (pi57 & w5557) | (pi57 & w8826) | (w5557 & w8826);
assign w5560 = ~w5557 & w8827;
assign w5561 = ~w5559 & ~w5560;
assign w5562 = (~w5376 & ~w5361) | (~w5376 & w8828) | (~w5361 & w8828);
assign w5563 = ~w5368 & ~w5562;
assign w5564 = ~w5562 & w7707;
assign w5565 = ~w5561 & ~w5563;
assign w5566 = ~w5564 & ~w5565;
assign w5567 = pi24 & w1132;
assign w5568 = pi23 & ~w1260;
assign w5569 = (pi51 & w5568) | (pi51 & w7708) | (w5568 & w7708);
assign w5570 = ~w5568 & w7709;
assign w5571 = ~w5569 & ~w5570;
assign w5572 = pi22 & w1393;
assign w5573 = pi21 & ~w2050;
assign w5574 = ~w2049 & w5573;
assign w5575 = ~w5572 & ~w5574;
assign w5576 = pi53 & ~w5575;
assign w5577 = ~pi53 & w5575;
assign w5578 = ~w5576 & ~w5577;
assign w5579 = pi20 & w1695;
assign w5580 = pi19 & ~w1865;
assign w5581 = ~w1864 & w5580;
assign w5582 = ~w5579 & ~w5581;
assign w5583 = pi55 & ~w5582;
assign w5584 = ~pi55 & w5582;
assign w5585 = ~w5583 & ~w5584;
assign w5586 = ~w5578 & ~w5585;
assign w5587 = w5578 & w5585;
assign w5588 = ~w5586 & ~w5587;
assign w5589 = w5571 & ~w5588;
assign w5590 = ~w5571 & w5588;
assign w5591 = ~w5589 & ~w5590;
assign w5592 = w5566 & ~w5591;
assign w5593 = ~w5566 & w5591;
assign w5594 = ~w5592 & ~w5593;
assign w5595 = ~w5556 & ~w5594;
assign w5596 = w5556 & w5594;
assign w5597 = ~w5595 & ~w5596;
assign w5598 = w5393 & ~w5416;
assign w5599 = ~w5393 & w5416;
assign w5600 = ~w5598 & ~w5599;
assign w5601 = ~w5431 & ~w5600;
assign w5602 = pi29 & ~w612;
assign w5603 = pi30 & w523;
assign w5604 = (pi45 & w5602) | (pi45 & w8829) | (w5602 & w8829);
assign w5605 = ~w5602 & w8830;
assign w5606 = ~w5604 & ~w5605;
assign w5607 = pi26 & w909;
assign w5608 = pi25 & ~w2273;
assign w5609 = ~w2272 & w5608;
assign w5610 = ~w5607 & ~w5609;
assign w5611 = pi49 & ~w5610;
assign w5612 = ~pi49 & w5610;
assign w5613 = ~w5611 & ~w5612;
assign w5614 = pi28 & w700;
assign w5615 = pi27 & ~w2099;
assign w5616 = ~w2098 & w5615;
assign w5617 = ~w5614 & ~w5616;
assign w5618 = pi47 & ~w5617;
assign w5619 = ~pi47 & w5617;
assign w5620 = ~w5618 & ~w5619;
assign w5621 = w5613 & w5620;
assign w5622 = ~w5613 & ~w5620;
assign w5623 = ~w5621 & ~w5622;
assign w5624 = w5606 & w5623;
assign w5625 = ~w5606 & ~w5623;
assign w5626 = ~w5624 & ~w5625;
assign w5627 = (~w5411 & ~w5413) | (~w5411 & w7710) | (~w5413 & w7710);
assign w5628 = w5626 & ~w5627;
assign w5629 = ~w5626 & w5627;
assign w5630 = ~w5628 & ~w5629;
assign w5631 = w5423 & ~w5630;
assign w5632 = ~w5423 & w5630;
assign w5633 = ~w5631 & ~w5632;
assign w5634 = ~w5601 & ~w5633;
assign w5635 = w5601 & w5633;
assign w5636 = ~w5634 & ~w5635;
assign w5637 = ~w5597 & w5636;
assign w5638 = w5597 & ~w5636;
assign w5639 = ~w5637 & ~w5638;
assign w5640 = w5550 & ~w5639;
assign w5641 = ~w5550 & w5639;
assign w5642 = ~w5640 & ~w5641;
assign w5643 = w5514 & ~w5642;
assign w5644 = ~w5514 & w5642;
assign w5645 = ~w5643 & ~w5644;
assign w5646 = ~w5505 & w5645;
assign w5647 = w5505 & ~w5645;
assign w5648 = ~w5646 & ~w5647;
assign w5649 = w5319 & w5497;
assign w5650 = w5320 & w8029;
assign w5651 = w4814 & w5650;
assign w5652 = (w5650 & w4817) | (w5650 & w7918) | (w4817 & w7918);
assign w5653 = ~w5318 & ~w5495;
assign w5654 = w4991 & w8831;
assign w5655 = (~w5317 & w5330) | (~w5317 & w7919) | (w5330 & w7919);
assign w5656 = ~w5654 & w5655;
assign w5657 = w4819 & w5321;
assign w5658 = w5656 & ~w5657;
assign w5659 = (~w5657 & w8832) | (~w5657 & w8833) | (w8832 & w8833);
assign w5660 = ~w5652 & w5659;
assign w5661 = (w5648 & w5651) | (w5648 & w7921) | (w5651 & w7921);
assign w5662 = ~w5651 & w8030;
assign w5663 = ~w5661 & ~w5662;
assign w5664 = (w5511 & ~w5514) | (w5511 & w7711) | (~w5514 & w7711);
assign w5665 = ~w5541 & ~w5544;
assign w5666 = ~w5548 & w5639;
assign w5667 = (w5665 & w5666) | (w5665 & w7712) | (w5666 & w7712);
assign w5668 = ~w5666 & w7713;
assign w5669 = ~w5667 & ~w5668;
assign w5670 = (~w5554 & ~w5556) | (~w5554 & w7714) | (~w5556 & w7714);
assign w5671 = (~w5532 & ~w5534) | (~w5532 & w8834) | (~w5534 & w8834);
assign w5672 = pi16 & ~w2588;
assign w5673 = pi17 & w2390;
assign w5674 = (pi59 & w5672) | (pi59 & w8835) | (w5672 & w8835);
assign w5675 = ~w5672 & w8836;
assign w5676 = ~w5674 & ~w5675;
assign w5677 = pi12 & ~w3404;
assign w5678 = pi13 & w3186;
assign w5679 = (pi63 & w5677) | (pi63 & w7922) | (w5677 & w7922);
assign w5680 = ~w5677 & w7923;
assign w5681 = ~w5679 & ~w5680;
assign w5682 = pi14 & ~w2981;
assign w5683 = pi15 & w2932;
assign w5684 = (pi61 & w5682) | (pi61 & w7924) | (w5682 & w7924);
assign w5685 = ~w5682 & w7925;
assign w5686 = ~w5684 & ~w5685;
assign w5687 = w5681 & w5686;
assign w5688 = ~w5681 & ~w5686;
assign w5689 = ~w5687 & ~w5688;
assign w5690 = w5676 & w5689;
assign w5691 = ~w5676 & ~w5689;
assign w5692 = ~w5690 & ~w5691;
assign w5693 = ~w5671 & w5692;
assign w5694 = w5671 & ~w5692;
assign w5695 = ~w5693 & ~w5694;
assign w5696 = w5538 & w5695;
assign w5697 = ~w5538 & ~w5695;
assign w5698 = ~w5696 & ~w5697;
assign w5699 = ~w5670 & w5698;
assign w5700 = w5670 & ~w5698;
assign w5701 = ~w5699 & ~w5700;
assign w5702 = (~w5634 & ~w5636) | (~w5634 & w8837) | (~w5636 & w8837);
assign w5703 = w5701 & w5702;
assign w5704 = ~w5701 & ~w5702;
assign w5705 = ~w5703 & ~w5704;
assign w5706 = (~w5621 & ~w5623) | (~w5621 & w8838) | (~w5623 & w8838);
assign w5707 = pi30 & ~w612;
assign w5708 = pi31 & ~w522;
assign w5709 = ~w521 & w5708;
assign w5710 = (pi45 & w5707) | (pi45 & w8839) | (w5707 & w8839);
assign w5711 = ~w5707 & w8840;
assign w5712 = ~w5710 & ~w5711;
assign w5713 = pi49 & w907;
assign w5714 = ~w2481 & ~w5713;
assign w5715 = pi26 & ~w5714;
assign w5716 = (pi49 & w5715) | (pi49 & w7715) | (w5715 & w7715);
assign w5717 = ~w5715 & w7716;
assign w5718 = ~w5716 & ~w5717;
assign w5719 = pi28 & ~w854;
assign w5720 = pi29 & w700;
assign w5721 = (pi47 & w5719) | (pi47 & w7717) | (w5719 & w7717);
assign w5722 = ~w5719 & w7718;
assign w5723 = ~w5721 & ~w5722;
assign w5724 = w5718 & w5723;
assign w5725 = ~w5718 & ~w5723;
assign w5726 = ~w5724 & ~w5725;
assign w5727 = w5712 & w5726;
assign w5728 = ~w5712 & ~w5726;
assign w5729 = ~w5727 & ~w5728;
assign w5730 = ~w5706 & w5729;
assign w5731 = w5706 & ~w5729;
assign w5732 = ~w5730 & ~w5731;
assign w5733 = w5423 & ~w5428;
assign w5734 = ~w5630 & w5733;
assign w5735 = w5429 & w5630;
assign w5736 = ~w5734 & ~w5735;
assign w5737 = w5732 & w5736;
assign w5738 = ~w5732 & ~w5736;
assign w5739 = ~w5737 & ~w5738;
assign w5740 = ~w5571 & ~w5587;
assign w5741 = pi19 & w2032;
assign w5742 = pi18 & ~w2206;
assign w5743 = (pi57 & w5742) | (pi57 & w7719) | (w5742 & w7719);
assign w5744 = ~w5742 & w7720;
assign w5745 = ~w5743 & ~w5744;
assign w5746 = ~w5586 & ~w5745;
assign w5747 = ~w5740 & w5746;
assign w5748 = w5571 & ~w5586;
assign w5749 = ~w5587 & w5745;
assign w5750 = ~w5748 & w5749;
assign w5751 = ~w5747 & ~w5750;
assign w5752 = pi21 & w1695;
assign w5753 = pi55 & w1693;
assign w5754 = ~w2428 & ~w5753;
assign w5755 = pi20 & ~w5754;
assign w5756 = (pi55 & w5755) | (pi55 & w7721) | (w5755 & w7721);
assign w5757 = ~w5755 & w7722;
assign w5758 = ~w5756 & ~w5757;
assign w5759 = pi25 & w1132;
assign w5760 = pi24 & ~w2419;
assign w5761 = ~w2418 & w5760;
assign w5762 = ~w5759 & ~w5761;
assign w5763 = pi51 & ~w5762;
assign w5764 = ~pi51 & w5762;
assign w5765 = ~w5763 & ~w5764;
assign w5766 = pi23 & w1393;
assign w5767 = pi22 & ~w2050;
assign w5768 = ~w2049 & w5767;
assign w5769 = ~w5766 & ~w5768;
assign w5770 = pi53 & ~w5769;
assign w5771 = ~pi53 & w5769;
assign w5772 = ~w5770 & ~w5771;
assign w5773 = ~w5765 & ~w5772;
assign w5774 = w5765 & w5772;
assign w5775 = ~w5773 & ~w5774;
assign w5776 = w5758 & ~w5775;
assign w5777 = ~w5758 & w5775;
assign w5778 = ~w5776 & ~w5777;
assign w5779 = ~w5751 & ~w5778;
assign w5780 = w5751 & w5778;
assign w5781 = ~w5779 & ~w5780;
assign w5782 = (~w5565 & ~w5591) | (~w5565 & w8841) | (~w5591 & w8841);
assign w5783 = ~w5781 & ~w5782;
assign w5784 = w5781 & w5782;
assign w5785 = ~w5783 & ~w5784;
assign w5786 = (~w5431 & ~w5626) | (~w5431 & w7926) | (~w5626 & w7926);
assign w5787 = ~w5629 & ~w5786;
assign w5788 = w5785 & ~w5787;
assign w5789 = ~w5785 & w5787;
assign w5790 = ~w5788 & ~w5789;
assign w5791 = w5739 & ~w5790;
assign w5792 = ~w5739 & w5790;
assign w5793 = ~w5791 & ~w5792;
assign w5794 = ~w5705 & w5793;
assign w5795 = w5705 & ~w5793;
assign w5796 = ~w5794 & ~w5795;
assign w5797 = w5669 & ~w5796;
assign w5798 = ~w5669 & w5796;
assign w5799 = ~w5797 & ~w5798;
assign w5800 = w5664 & w5799;
assign w5801 = ~w5664 & ~w5799;
assign w5802 = ~w5800 & ~w5801;
assign w5803 = w5661 & w5802;
assign w5804 = w5647 & ~w5802;
assign w5805 = ~w5647 & w5802;
assign w5806 = ~w5804 & ~w5805;
assign w5807 = ~w5661 & w5806;
assign w5808 = ~w5803 & ~w5807;
assign w5809 = ~w5703 & ~w5793;
assign w5810 = ~w5696 & ~w5699;
assign w5811 = (~w5810 & w5702) | (~w5810 & w7723) | (w5702 & w7723);
assign w5812 = ~w5809 & w5811;
assign w5813 = ~w5704 & w5793;
assign w5814 = (w5810 & ~w5702) | (w5810 & w7724) | (~w5702 & w7724);
assign w5815 = ~w5813 & w5814;
assign w5816 = ~w5812 & ~w5815;
assign w5817 = (~w5687 & ~w5689) | (~w5687 & w8842) | (~w5689 & w8842);
assign w5818 = pi17 & ~w2588;
assign w5819 = pi18 & w2390;
assign w5820 = (pi59 & w5818) | (pi59 & w8843) | (w5818 & w8843);
assign w5821 = ~w5818 & w8844;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = pi13 & ~w3404;
assign w5824 = pi14 & w3186;
assign w5825 = (pi63 & w5823) | (pi63 & w7927) | (w5823 & w7927);
assign w5826 = ~w5823 & w7928;
assign w5827 = ~w5825 & ~w5826;
assign w5828 = pi15 & ~w2981;
assign w5829 = pi16 & w2932;
assign w5830 = (pi61 & w5828) | (pi61 & w7929) | (w5828 & w7929);
assign w5831 = ~w5828 & w7930;
assign w5832 = ~w5830 & ~w5831;
assign w5833 = w5827 & w5832;
assign w5834 = ~w5827 & ~w5832;
assign w5835 = ~w5833 & ~w5834;
assign w5836 = w5822 & w5835;
assign w5837 = ~w5822 & ~w5835;
assign w5838 = ~w5836 & ~w5837;
assign w5839 = w5817 & ~w5838;
assign w5840 = ~w5817 & w5838;
assign w5841 = ~w5839 & ~w5840;
assign w5842 = w5693 & w5841;
assign w5843 = ~w5693 & ~w5841;
assign w5844 = ~w5842 & ~w5843;
assign w5845 = (~w5783 & ~w5785) | (~w5783 & w7725) | (~w5785 & w7725);
assign w5846 = ~w5844 & ~w5845;
assign w5847 = w5844 & w5845;
assign w5848 = ~w5846 & ~w5847;
assign w5849 = w5745 & ~w5750;
assign w5850 = ~w5779 & ~w5849;
assign w5851 = pi19 & ~w2206;
assign w5852 = pi20 & w2032;
assign w5853 = (pi57 & w5851) | (pi57 & w7931) | (w5851 & w7931);
assign w5854 = ~w5851 & w7932;
assign w5855 = ~w5853 & ~w5854;
assign w5856 = ~w5758 & ~w5774;
assign w5857 = ~w5856 & w7726;
assign w5858 = (~w5855 & w5856) | (~w5855 & w7727) | (w5856 & w7727);
assign w5859 = ~w5857 & ~w5858;
assign w5860 = pi26 & w1132;
assign w5861 = pi25 & ~w1260;
assign w5862 = (pi51 & w5861) | (pi51 & w7728) | (w5861 & w7728);
assign w5863 = ~w5861 & w7729;
assign w5864 = ~w5862 & ~w5863;
assign w5865 = pi24 & w1393;
assign w5866 = pi23 & ~w2050;
assign w5867 = ~w2049 & w5866;
assign w5868 = ~w5865 & ~w5867;
assign w5869 = pi53 & ~w5868;
assign w5870 = ~pi53 & w5868;
assign w5871 = ~w5869 & ~w5870;
assign w5872 = pi22 & w1695;
assign w5873 = pi21 & ~w1865;
assign w5874 = ~w1864 & w5873;
assign w5875 = ~w5872 & ~w5874;
assign w5876 = pi55 & ~w5875;
assign w5877 = ~pi55 & w5875;
assign w5878 = ~w5876 & ~w5877;
assign w5879 = ~w5871 & ~w5878;
assign w5880 = w5871 & w5878;
assign w5881 = ~w5879 & ~w5880;
assign w5882 = w5864 & ~w5881;
assign w5883 = ~w5864 & w5881;
assign w5884 = ~w5882 & ~w5883;
assign w5885 = w5859 & w5884;
assign w5886 = ~w5859 & ~w5884;
assign w5887 = ~w5885 & ~w5886;
assign w5888 = ~w5850 & ~w5887;
assign w5889 = w5850 & w5887;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = (~w5724 & ~w5726) | (~w5724 & w7933) | (~w5726 & w7933);
assign w5892 = pi27 & ~w5714;
assign w5893 = (pi49 & w5892) | (pi49 & w7730) | (w5892 & w7730);
assign w5894 = ~w5892 & w7731;
assign w5895 = ~w5893 & ~w5894;
assign w5896 = pi29 & ~w854;
assign w5897 = (pi47 & w5896) | (pi47 & w7732) | (w5896 & w7732);
assign w5898 = ~w5896 & w7733;
assign w5899 = ~w5897 & ~w5898;
assign w5900 = w5895 & w5899;
assign w5901 = ~w5895 & ~w5899;
assign w5902 = ~w5900 & ~w5901;
assign w5903 = (pi45 & w522) | (pi45 & w8845) | (w522 & w8845);
assign w5904 = pi31 & ~pi45;
assign w5905 = ~w521 & w5904;
assign w5906 = ~w5903 & ~w5905;
assign w5907 = ~w5902 & ~w5906;
assign w5908 = w5902 & w5906;
assign w5909 = ~w5907 & ~w5908;
assign w5910 = ~w5891 & w5909;
assign w5911 = w5891 & ~w5909;
assign w5912 = ~w5910 & ~w5911;
assign w5913 = ~w5731 & w5912;
assign w5914 = w5731 & ~w5912;
assign w5915 = ~w5913 & ~w5914;
assign w5916 = w5890 & ~w5915;
assign w5917 = ~w5890 & w5915;
assign w5918 = ~w5916 & ~w5917;
assign w5919 = ~w5791 & w7734;
assign w5920 = (~w5918 & w5791) | (~w5918 & w7735) | (w5791 & w7735);
assign w5921 = ~w5919 & ~w5920;
assign w5922 = w5848 & ~w5921;
assign w5923 = ~w5848 & w5921;
assign w5924 = ~w5922 & ~w5923;
assign w5925 = w5816 & ~w5924;
assign w5926 = ~w5816 & w5924;
assign w5927 = ~w5925 & ~w5926;
assign w5928 = (~w5667 & ~w5796) | (~w5667 & w7736) | (~w5796 & w7736);
assign w5929 = ~w5927 & ~w5928;
assign w5930 = w5927 & w5928;
assign w5931 = ~w5929 & ~w5930;
assign w5932 = ~w5646 & w5653;
assign w5933 = ~w5649 & w5932;
assign w5934 = ~w5496 & ~w5647;
assign w5935 = ~w5646 & ~w5934;
assign w5936 = (~w5800 & w5934) | (~w5800 & w7737) | (w5934 & w7737);
assign w5937 = ~w5933 & w5936;
assign w5938 = (~w5801 & w5933) | (~w5801 & w8846) | (w5933 & w8846);
assign w5939 = w5648 & ~w5800;
assign w5940 = w5649 & w5939;
assign w5941 = w5331 & w5940;
assign w5942 = ~w5938 & ~w5941;
assign w5943 = ~w5801 & ~w5942;
assign w5944 = ~w4994 & ~w5943;
assign w5945 = w5648 & w5802;
assign w5946 = w5649 & w5945;
assign w5947 = w5945 & w7738;
assign w5948 = (~w5947 & w5942) | (~w5947 & w8031) | (w5942 & w8031);
assign w5949 = (~w5948 & w5000) | (~w5948 & w7934) | (w5000 & w7934);
assign w5950 = w5931 & ~w5949;
assign w5951 = ~w5931 & w5949;
assign w5952 = ~w5950 & ~w5951;
assign w5953 = (~w5812 & ~w5816) | (~w5812 & w7739) | (~w5816 & w7739);
assign w5954 = w5842 & w5845;
assign w5955 = ~w5919 & w5954;
assign w5956 = (~w5842 & ~w5845) | (~w5842 & w7935) | (~w5845 & w7935);
assign w5957 = w5920 & ~w5956;
assign w5958 = ~w5955 & ~w5957;
assign w5959 = (~w5846 & w5791) | (~w5846 & w7740) | (w5791 & w7740);
assign w5960 = w5918 & w5956;
assign w5961 = ~w5959 & w5960;
assign w5962 = w5843 & ~w5845;
assign w5963 = ~w5791 & w7936;
assign w5964 = ~w5961 & ~w5963;
assign w5965 = w5958 & w5964;
assign w5966 = (~w5833 & ~w5835) | (~w5833 & w8847) | (~w5835 & w8847);
assign w5967 = pi18 & ~w2588;
assign w5968 = pi19 & w2390;
assign w5969 = (pi59 & w5967) | (pi59 & w8848) | (w5967 & w8848);
assign w5970 = ~w5967 & w8849;
assign w5971 = ~w5969 & ~w5970;
assign w5972 = pi14 & ~w3404;
assign w5973 = pi15 & w3186;
assign w5974 = (pi63 & w5972) | (pi63 & w7741) | (w5972 & w7741);
assign w5975 = ~w5972 & w7742;
assign w5976 = ~w5974 & ~w5975;
assign w5977 = pi16 & ~w2981;
assign w5978 = pi17 & w2932;
assign w5979 = (pi61 & w5977) | (pi61 & w7743) | (w5977 & w7743);
assign w5980 = ~w5977 & w7744;
assign w5981 = ~w5979 & ~w5980;
assign w5982 = w5976 & w5981;
assign w5983 = ~w5976 & ~w5981;
assign w5984 = ~w5982 & ~w5983;
assign w5985 = w5971 & w5984;
assign w5986 = ~w5971 & ~w5984;
assign w5987 = ~w5985 & ~w5986;
assign w5988 = ~w5966 & w5987;
assign w5989 = w5966 & ~w5987;
assign w5990 = ~w5988 & ~w5989;
assign w5991 = w5840 & w5990;
assign w5992 = ~w5840 & ~w5990;
assign w5993 = ~w5991 & ~w5992;
assign w5994 = ~w5730 & ~w5888;
assign w5995 = ~w5889 & ~w5994;
assign w5996 = w5993 & w5995;
assign w5997 = ~w5993 & ~w5995;
assign w5998 = ~w5996 & ~w5997;
assign w5999 = ~w5864 & ~w5880;
assign w6000 = pi21 & w2032;
assign w6001 = pi20 & ~w2206;
assign w6002 = (pi57 & w6001) | (pi57 & w7745) | (w6001 & w7745);
assign w6003 = ~w6001 & w7746;
assign w6004 = ~w6002 & ~w6003;
assign w6005 = ~w5879 & ~w6004;
assign w6006 = ~w5999 & w6005;
assign w6007 = w5864 & ~w5879;
assign w6008 = ~w5880 & w6004;
assign w6009 = ~w6007 & w6008;
assign w6010 = ~w6006 & ~w6009;
assign w6011 = pi27 & w1132;
assign w6012 = pi26 & ~w1260;
assign w6013 = (pi51 & w6012) | (pi51 & w7747) | (w6012 & w7747);
assign w6014 = ~w6012 & w7748;
assign w6015 = ~w6013 & ~w6014;
assign w6016 = pi25 & w1393;
assign w6017 = pi24 & ~w2050;
assign w6018 = ~w2049 & w6017;
assign w6019 = ~w6016 & ~w6018;
assign w6020 = pi53 & ~w6019;
assign w6021 = ~pi53 & w6019;
assign w6022 = ~w6020 & ~w6021;
assign w6023 = pi23 & w1695;
assign w6024 = pi22 & ~w1865;
assign w6025 = ~w1864 & w6024;
assign w6026 = ~w6023 & ~w6025;
assign w6027 = pi55 & ~w6026;
assign w6028 = ~pi55 & w6026;
assign w6029 = ~w6027 & ~w6028;
assign w6030 = ~w6022 & ~w6029;
assign w6031 = w6022 & w6029;
assign w6032 = ~w6030 & ~w6031;
assign w6033 = w6015 & ~w6032;
assign w6034 = ~w6015 & w6032;
assign w6035 = ~w6033 & ~w6034;
assign w6036 = ~w6010 & ~w6035;
assign w6037 = w6010 & w6035;
assign w6038 = ~w6036 & ~w6037;
assign w6039 = (~w5857 & w5884) | (~w5857 & w7749) | (w5884 & w7749);
assign w6040 = ~w6038 & w6039;
assign w6041 = w6038 & ~w6039;
assign w6042 = ~w6040 & ~w6041;
assign w6043 = (~w5900 & ~w5902) | (~w5900 & w7937) | (~w5902 & w7937);
assign w6044 = pi28 & ~w5714;
assign w6045 = pi29 & w909;
assign w6046 = (pi49 & w6044) | (pi49 & w8850) | (w6044 & w8850);
assign w6047 = ~w6044 & w8851;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = pi30 & ~w854;
assign w6050 = pi31 & ~w699;
assign w6051 = ~w698 & w6050;
assign w6052 = (pi47 & w6049) | (pi47 & w8852) | (w6049 & w8852);
assign w6053 = ~w6049 & w8853;
assign w6054 = ~w6052 & ~w6053;
assign w6055 = w6048 & w6054;
assign w6056 = ~w6048 & ~w6054;
assign w6057 = ~w6055 & ~w6056;
assign w6058 = ~w6043 & ~w6057;
assign w6059 = w6043 & w6057;
assign w6060 = ~w6058 & ~w6059;
assign w6061 = ~w5910 & w6060;
assign w6062 = w5910 & ~w6060;
assign w6063 = ~w6061 & ~w6062;
assign w6064 = w6042 & w6063;
assign w6065 = ~w6042 & ~w6063;
assign w6066 = ~w6064 & ~w6065;
assign w6067 = ~w5890 & w5913;
assign w6068 = (~w5730 & w5912) | (~w5730 & w5732) | (w5912 & w5732);
assign w6069 = w5890 & w6068;
assign w6070 = ~w6067 & ~w6069;
assign w6071 = ~w6066 & ~w6070;
assign w6072 = w6066 & w6070;
assign w6073 = ~w6071 & ~w6072;
assign w6074 = w5998 & ~w6073;
assign w6075 = ~w5998 & w6073;
assign w6076 = ~w6074 & ~w6075;
assign w6077 = ~w5965 & w6076;
assign w6078 = w5965 & ~w6076;
assign w6079 = ~w6077 & ~w6078;
assign w6080 = w5953 & ~w6079;
assign w6081 = ~w5953 & w6079;
assign w6082 = ~w6080 & ~w6081;
assign w6083 = w5930 & ~w6082;
assign w6084 = ~w5930 & w6082;
assign w6085 = ~w6083 & ~w6084;
assign w6086 = w5931 & w6082;
assign w6087 = (~w6086 & ~w6085) | (~w6086 & w8854) | (~w6085 & w8854);
assign w6088 = w5949 & ~w6087;
assign w6089 = ~w5949 & w6085;
assign w6090 = ~w6088 & ~w6089;
assign w6091 = ~w5331 & ~w5938;
assign w6092 = (w6091 & w5333) | (w6091 & w8855) | (w5333 & w8855);
assign w6093 = (w6086 & w5938) | (w6086 & w8032) | (w5938 & w8032);
assign w6094 = (w5958 & ~w5965) | (w5958 & w7938) | (~w5965 & w7938);
assign w6095 = (~w5991 & ~w5995) | (~w5991 & w8856) | (~w5995 & w8856);
assign w6096 = w5998 & ~w6072;
assign w6097 = ~w6096 & w7939;
assign w6098 = (~w6095 & w6096) | (~w6095 & w7940) | (w6096 & w7940);
assign w6099 = ~w6097 & ~w6098;
assign w6100 = w6042 & w6061;
assign w6101 = w5910 & w6060;
assign w6102 = ~w6042 & w6101;
assign w6103 = ~w6100 & ~w6102;
assign w6104 = w6004 & ~w6009;
assign w6105 = ~w6036 & ~w6104;
assign w6106 = ~w6015 & ~w6031;
assign w6107 = pi22 & w2032;
assign w6108 = pi21 & ~w2206;
assign w6109 = (pi57 & w6108) | (pi57 & w7750) | (w6108 & w7750);
assign w6110 = ~w6108 & w7751;
assign w6111 = ~w6109 & ~w6110;
assign w6112 = ~w6030 & ~w6111;
assign w6113 = ~w6106 & w6112;
assign w6114 = w6015 & ~w6030;
assign w6115 = ~w6031 & w6111;
assign w6116 = ~w6114 & w6115;
assign w6117 = ~w6113 & ~w6116;
assign w6118 = pi24 & w1695;
assign w6119 = pi23 & ~w5754;
assign w6120 = (pi55 & w6119) | (pi55 & w7752) | (w6119 & w7752);
assign w6121 = ~w6119 & w7753;
assign w6122 = ~w6120 & ~w6121;
assign w6123 = pi28 & w1132;
assign w6124 = pi27 & ~w2419;
assign w6125 = ~w2418 & w6124;
assign w6126 = ~w6123 & ~w6125;
assign w6127 = pi51 & ~w6126;
assign w6128 = ~pi51 & w6126;
assign w6129 = ~w6127 & ~w6128;
assign w6130 = pi26 & w1393;
assign w6131 = pi25 & ~w2050;
assign w6132 = ~w2049 & w6131;
assign w6133 = ~w6130 & ~w6132;
assign w6134 = pi53 & ~w6133;
assign w6135 = ~pi53 & w6133;
assign w6136 = ~w6134 & ~w6135;
assign w6137 = ~w6129 & ~w6136;
assign w6138 = w6129 & w6136;
assign w6139 = ~w6137 & ~w6138;
assign w6140 = w6122 & ~w6139;
assign w6141 = ~w6122 & w6139;
assign w6142 = ~w6140 & ~w6141;
assign w6143 = ~w6117 & ~w6142;
assign w6144 = w6117 & w6142;
assign w6145 = ~w6143 & ~w6144;
assign w6146 = w6105 & ~w6145;
assign w6147 = ~w6105 & w6145;
assign w6148 = ~w6146 & ~w6147;
assign w6149 = pi29 & ~w5714;
assign w6150 = pi30 & w909;
assign w6151 = (pi49 & w6149) | (pi49 & w7754) | (w6149 & w7754);
assign w6152 = ~w6149 & w7755;
assign w6153 = ~w6151 & ~w6152;
assign w6154 = (pi47 & w699) | (pi47 & w8857) | (w699 & w8857);
assign w6155 = pi31 & ~pi47;
assign w6156 = ~w698 & w6155;
assign w6157 = ~w6154 & ~w6156;
assign w6158 = w6153 & w6157;
assign w6159 = ~w6153 & ~w6157;
assign w6160 = ~w6158 & ~w6159;
assign w6161 = w6056 & ~w6160;
assign w6162 = ~w6056 & w6160;
assign w6163 = ~w6161 & ~w6162;
assign w6164 = w6058 & w6163;
assign w6165 = ~w6058 & ~w6163;
assign w6166 = ~w6164 & ~w6165;
assign w6167 = w6148 & w6166;
assign w6168 = ~w6148 & ~w6166;
assign w6169 = ~w6167 & ~w6168;
assign w6170 = w6103 & ~w6169;
assign w6171 = ~w6103 & w6169;
assign w6172 = ~w6170 & ~w6171;
assign w6173 = (~w5982 & ~w5984) | (~w5982 & w8858) | (~w5984 & w8858);
assign w6174 = pi19 & ~w2588;
assign w6175 = pi20 & w2390;
assign w6176 = (pi59 & w6174) | (pi59 & w8859) | (w6174 & w8859);
assign w6177 = ~w6174 & w8860;
assign w6178 = ~w6176 & ~w6177;
assign w6179 = pi15 & ~w3404;
assign w6180 = pi16 & w3186;
assign w6181 = (pi63 & w6179) | (pi63 & w7756) | (w6179 & w7756);
assign w6182 = ~w6179 & w7757;
assign w6183 = ~w6181 & ~w6182;
assign w6184 = pi17 & ~w2981;
assign w6185 = pi18 & w2932;
assign w6186 = (pi61 & w6184) | (pi61 & w7758) | (w6184 & w7758);
assign w6187 = ~w6184 & w7759;
assign w6188 = ~w6186 & ~w6187;
assign w6189 = w6183 & w6188;
assign w6190 = ~w6183 & ~w6188;
assign w6191 = ~w6189 & ~w6190;
assign w6192 = w6178 & w6191;
assign w6193 = ~w6178 & ~w6191;
assign w6194 = ~w6192 & ~w6193;
assign w6195 = w6173 & ~w6194;
assign w6196 = ~w6173 & w6194;
assign w6197 = ~w6195 & ~w6196;
assign w6198 = w5988 & w6197;
assign w6199 = ~w5988 & ~w6197;
assign w6200 = ~w6198 & ~w6199;
assign w6201 = (w5910 & w6038) | (w5910 & w7760) | (w6038 & w7760);
assign w6202 = ~w6041 & ~w6201;
assign w6203 = w6200 & ~w6202;
assign w6204 = ~w6200 & w6202;
assign w6205 = ~w6203 & ~w6204;
assign w6206 = ~w6172 & w6205;
assign w6207 = w6172 & ~w6205;
assign w6208 = ~w6206 & ~w6207;
assign w6209 = w6099 & w6208;
assign w6210 = ~w6099 & ~w6208;
assign w6211 = ~w6209 & ~w6210;
assign w6212 = ~w6094 & ~w6211;
assign w6213 = w6094 & w6211;
assign w6214 = ~w6212 & ~w6213;
assign w6215 = (~w6080 & w5930) | (~w6080 & w7761) | (w5930 & w7761);
assign w6216 = ~w6214 & ~w6215;
assign w6217 = (w5329 & w8058) | (w5329 & w8059) | (w8058 & w8059);
assign w6218 = w6093 & w6214;
assign w6219 = (w6218 & ~w5329) | (w6218 & w7941) | (~w5329 & w7941);
assign w6220 = ~w6080 & w9086;
assign w6221 = ~w6219 & ~w6220;
assign w6222 = ~w6217 & w6221;
assign w6223 = ~w6198 & ~w6203;
assign w6224 = ~w6170 & w6205;
assign w6225 = ~w6224 & w7762;
assign w6226 = (~w6223 & w6224) | (~w6223 & w7763) | (w6224 & w7763);
assign w6227 = ~w6225 & ~w6226;
assign w6228 = ~w6148 & w6164;
assign w6229 = ~w6058 & w6163;
assign w6230 = w6148 & w6229;
assign w6231 = ~w6228 & ~w6230;
assign w6232 = (~w6189 & ~w6191) | (~w6189 & w8862) | (~w6191 & w8862);
assign w6233 = pi20 & ~w2588;
assign w6234 = pi21 & w2390;
assign w6235 = (pi59 & w6233) | (pi59 & w8863) | (w6233 & w8863);
assign w6236 = ~w6233 & w8864;
assign w6237 = ~w6235 & ~w6236;
assign w6238 = pi16 & ~w3404;
assign w6239 = pi17 & w3186;
assign w6240 = (pi63 & w6238) | (pi63 & w7764) | (w6238 & w7764);
assign w6241 = ~w6238 & w7765;
assign w6242 = ~w6240 & ~w6241;
assign w6243 = pi18 & ~w2981;
assign w6244 = pi19 & w2932;
assign w6245 = (pi61 & w6243) | (pi61 & w7766) | (w6243 & w7766);
assign w6246 = ~w6243 & w7767;
assign w6247 = ~w6245 & ~w6246;
assign w6248 = w6242 & w6247;
assign w6249 = ~w6242 & ~w6247;
assign w6250 = ~w6248 & ~w6249;
assign w6251 = w6237 & w6250;
assign w6252 = ~w6237 & ~w6250;
assign w6253 = ~w6251 & ~w6252;
assign w6254 = ~w6232 & w6253;
assign w6255 = w6232 & ~w6253;
assign w6256 = ~w6254 & ~w6255;
assign w6257 = w6196 & w6256;
assign w6258 = ~w6196 & ~w6256;
assign w6259 = ~w6257 & ~w6258;
assign w6260 = ~w6058 & ~w6147;
assign w6261 = ~w6146 & ~w6260;
assign w6262 = w6259 & w6261;
assign w6263 = ~w6259 & ~w6261;
assign w6264 = ~w6262 & ~w6263;
assign w6265 = pi22 & ~w2206;
assign w6266 = pi23 & w2032;
assign w6267 = (pi57 & w6265) | (pi57 & w8865) | (w6265 & w8865);
assign w6268 = ~w6265 & w8866;
assign w6269 = ~w6267 & ~w6268;
assign w6270 = ~w6122 & ~w6138;
assign w6271 = ~w6270 & w7768;
assign w6272 = (~w6269 & w6270) | (~w6269 & w7769) | (w6270 & w7769);
assign w6273 = ~w6271 & ~w6272;
assign w6274 = pi29 & w1132;
assign w6275 = pi28 & ~w1260;
assign w6276 = (pi51 & w6275) | (pi51 & w7770) | (w6275 & w7770);
assign w6277 = ~w6275 & w7771;
assign w6278 = ~w6276 & ~w6277;
assign w6279 = pi27 & w1393;
assign w6280 = pi26 & ~w2050;
assign w6281 = ~w2049 & w6280;
assign w6282 = ~w6279 & ~w6281;
assign w6283 = pi53 & ~w6282;
assign w6284 = ~pi53 & w6282;
assign w6285 = ~w6283 & ~w6284;
assign w6286 = pi25 & w1695;
assign w6287 = pi24 & ~w1865;
assign w6288 = ~w1864 & w6287;
assign w6289 = ~w6286 & ~w6288;
assign w6290 = pi55 & ~w6289;
assign w6291 = ~pi55 & w6289;
assign w6292 = ~w6290 & ~w6291;
assign w6293 = ~w6285 & ~w6292;
assign w6294 = w6285 & w6292;
assign w6295 = ~w6293 & ~w6294;
assign w6296 = w6278 & ~w6295;
assign w6297 = ~w6278 & w6295;
assign w6298 = ~w6296 & ~w6297;
assign w6299 = w6273 & w6298;
assign w6300 = ~w6273 & ~w6298;
assign w6301 = ~w6299 & ~w6300;
assign w6302 = w6111 & ~w6116;
assign w6303 = ~w6143 & ~w6302;
assign w6304 = pi30 & ~w5714;
assign w6305 = pi31 & ~w908;
assign w6306 = ~w907 & w6305;
assign w6307 = (pi49 & w6304) | (pi49 & w8867) | (w6304 & w8867);
assign w6308 = ~w6304 & w8868;
assign w6309 = ~w6307 & ~w6308;
assign w6310 = w6160 & w8869;
assign w6311 = w6158 & ~w6309;
assign w6312 = ~w6158 & w6309;
assign w6313 = ~w6311 & ~w6312;
assign w6314 = ~w6162 & ~w6313;
assign w6315 = ~w6310 & ~w6314;
assign w6316 = w6303 & ~w6315;
assign w6317 = ~w6303 & w6315;
assign w6318 = ~w6316 & ~w6317;
assign w6319 = w6301 & w6318;
assign w6320 = ~w6301 & ~w6318;
assign w6321 = ~w6319 & ~w6320;
assign w6322 = w6264 & ~w6321;
assign w6323 = ~w6264 & w6321;
assign w6324 = ~w6322 & ~w6323;
assign w6325 = w6231 & ~w6324;
assign w6326 = ~w6231 & ~w6321;
assign w6327 = ~w6264 & w6326;
assign w6328 = ~w6231 & w6321;
assign w6329 = w6264 & w6328;
assign w6330 = ~w6327 & ~w6329;
assign w6331 = ~w6325 & w6330;
assign w6332 = w6227 & ~w6331;
assign w6333 = ~w6227 & w6331;
assign w6334 = ~w6332 & ~w6333;
assign w6335 = (~w6098 & w6208) | (~w6098 & w8870) | (w6208 & w8870);
assign w6336 = w6334 & w6335;
assign w6337 = ~w6334 & ~w6335;
assign w6338 = ~w6336 & ~w6337;
assign w6339 = (~w6212 & ~w6215) | (~w6212 & w8033) | (~w6215 & w8033);
assign w6340 = ~w5334 & w7942;
assign w6341 = (w5329 & w8034) | (w5329 & w8035) | (w8034 & w8035);
assign w6342 = (w7944 & ~w5329) | (w7944 & w8036) | (~w5329 & w8036);
assign w6343 = ~w6341 & ~w6342;
assign w6344 = (~w6257 & ~w6261) | (~w6257 & w8871) | (~w6261 & w8871);
assign w6345 = (w6344 & ~w6264) | (w6344 & w8872) | (~w6264 & w8872);
assign w6346 = w6330 & w6345;
assign w6347 = (w6231 & ~w6264) | (w6231 & w7772) | (~w6264 & w7772);
assign w6348 = (~w6344 & w6264) | (~w6344 & w8873) | (w6264 & w8873);
assign w6349 = ~w6347 & w6348;
assign w6350 = ~w6346 & ~w6349;
assign w6351 = (~w6248 & ~w6250) | (~w6248 & w8874) | (~w6250 & w8874);
assign w6352 = pi21 & ~w2588;
assign w6353 = pi22 & w2390;
assign w6354 = (pi59 & w6352) | (pi59 & w8875) | (w6352 & w8875);
assign w6355 = ~w6352 & w8876;
assign w6356 = ~w6354 & ~w6355;
assign w6357 = pi17 & ~w3404;
assign w6358 = pi18 & w3186;
assign w6359 = (pi63 & w6357) | (pi63 & w7773) | (w6357 & w7773);
assign w6360 = ~w6357 & w7774;
assign w6361 = ~w6359 & ~w6360;
assign w6362 = pi19 & ~w2981;
assign w6363 = pi20 & w2932;
assign w6364 = (pi61 & w6362) | (pi61 & w7775) | (w6362 & w7775);
assign w6365 = ~w6362 & w7776;
assign w6366 = ~w6364 & ~w6365;
assign w6367 = w6361 & w6366;
assign w6368 = ~w6361 & ~w6366;
assign w6369 = ~w6367 & ~w6368;
assign w6370 = w6356 & w6369;
assign w6371 = ~w6356 & ~w6369;
assign w6372 = ~w6370 & ~w6371;
assign w6373 = ~w6351 & w6372;
assign w6374 = w6351 & ~w6372;
assign w6375 = ~w6373 & ~w6374;
assign w6376 = w6254 & w6375;
assign w6377 = ~w6254 & ~w6375;
assign w6378 = ~w6376 & ~w6377;
assign w6379 = (w6162 & w6143) | (w6162 & w8877) | (w6143 & w8877);
assign w6380 = ~w6143 & w7777;
assign w6381 = ~w6301 & ~w6380;
assign w6382 = ~w6379 & ~w6381;
assign w6383 = ~w6378 & w6382;
assign w6384 = w6378 & ~w6382;
assign w6385 = ~w6383 & ~w6384;
assign w6386 = w6313 & w6321;
assign w6387 = ~w6385 & ~w6386;
assign w6388 = w6385 & w6386;
assign w6389 = ~w6387 & ~w6388;
assign w6390 = ~w6278 & ~w6294;
assign w6391 = pi24 & w2032;
assign w6392 = pi23 & ~w2206;
assign w6393 = (pi57 & w6392) | (pi57 & w7778) | (w6392 & w7778);
assign w6394 = ~w6392 & w7779;
assign w6395 = ~w6393 & ~w6394;
assign w6396 = ~w6293 & ~w6395;
assign w6397 = ~w6390 & w6396;
assign w6398 = w6278 & ~w6293;
assign w6399 = ~w6294 & w6395;
assign w6400 = ~w6398 & w6399;
assign w6401 = ~w6397 & ~w6400;
assign w6402 = pi30 & w1132;
assign w6403 = pi29 & ~w1260;
assign w6404 = (pi51 & w6403) | (pi51 & w7780) | (w6403 & w7780);
assign w6405 = ~w6403 & w7781;
assign w6406 = ~w6404 & ~w6405;
assign w6407 = pi28 & w1393;
assign w6408 = pi27 & ~w2050;
assign w6409 = ~w2049 & w6408;
assign w6410 = ~w6407 & ~w6409;
assign w6411 = pi53 & ~w6410;
assign w6412 = ~pi53 & w6410;
assign w6413 = ~w6411 & ~w6412;
assign w6414 = pi26 & w1695;
assign w6415 = pi25 & ~w1865;
assign w6416 = ~w1864 & w6415;
assign w6417 = ~w6414 & ~w6416;
assign w6418 = pi55 & ~w6417;
assign w6419 = ~pi55 & w6417;
assign w6420 = ~w6418 & ~w6419;
assign w6421 = ~w6413 & ~w6420;
assign w6422 = w6413 & w6420;
assign w6423 = ~w6421 & ~w6422;
assign w6424 = w6406 & ~w6423;
assign w6425 = ~w6406 & w6423;
assign w6426 = ~w6424 & ~w6425;
assign w6427 = ~w6401 & ~w6426;
assign w6428 = w6401 & w6426;
assign w6429 = ~w6427 & ~w6428;
assign w6430 = (~w6271 & w6298) | (~w6271 & w7782) | (w6298 & w7782);
assign w6431 = w6429 & ~w6430;
assign w6432 = ~w6429 & w6430;
assign w6433 = ~w6431 & ~w6432;
assign w6434 = (pi49 & w908) | (pi49 & w8878) | (w908 & w8878);
assign w6435 = pi31 & ~pi49;
assign w6436 = ~w907 & w6435;
assign w6437 = ~w6434 & ~w6436;
assign w6438 = w6309 & w6437;
assign w6439 = ~w6309 & ~w6437;
assign w6440 = ~w6438 & ~w6439;
assign w6441 = ~w6311 & w6440;
assign w6442 = w6433 & w6441;
assign w6443 = w6158 & w8879;
assign w6444 = ~w6433 & w6443;
assign w6445 = ~w6442 & ~w6444;
assign w6446 = (~w6311 & ~w6429) | (~w6311 & w7783) | (~w6429 & w7783);
assign w6447 = ~w6432 & w6446;
assign w6448 = (~w6440 & w6433) | (~w6440 & w7784) | (w6433 & w7784);
assign w6449 = ~w6447 & w6448;
assign w6450 = w6445 & ~w6449;
assign w6451 = ~w6389 & w6450;
assign w6452 = w6389 & ~w6450;
assign w6453 = ~w6451 & ~w6452;
assign w6454 = ~w6350 & w6453;
assign w6455 = w6350 & ~w6453;
assign w6456 = ~w6454 & ~w6455;
assign w6457 = (~w6225 & w6331) | (~w6225 & w7785) | (w6331 & w7785);
assign w6458 = ~w6456 & ~w6457;
assign w6459 = w6456 & w6457;
assign w6460 = ~w6458 & ~w6459;
assign w6461 = ~w5801 & w6214;
assign w6462 = w6086 & w6461;
assign w6463 = w6086 & w7945;
assign w6464 = w5648 & w6463;
assign w6465 = w5650 & w6464;
assign w6466 = w4813 & w6465;
assign w6467 = (w6466 & w3602) | (w6466 & w8037) | (w3602 & w8037);
assign w6468 = (w6465 & w4817) | (w6465 & w8038) | (w4817 & w8038);
assign w6469 = (~w8037 & w9074) | (~w8037 & w9075) | (w9074 & w9075);
assign w6470 = w6463 & w8880;
assign w6471 = w6086 & w7786;
assign w6472 = ~w6471 & w8039;
assign w6473 = w5935 & w6463;
assign w6474 = w6472 & ~w6473;
assign w6475 = (w6474 & w5658) | (w6474 & w8040) | (w5658 & w8040);
assign w6476 = ~w6467 & w7787;
assign w6477 = (w6460 & w6476) | (w6460 & w7946) | (w6476 & w7946);
assign w6478 = ~w6476 & w7947;
assign w6479 = ~w6477 & ~w6478;
assign w6480 = ~w6349 & ~w6455;
assign w6481 = ~w6376 & ~w6384;
assign w6482 = ~w6388 & ~w6450;
assign w6483 = (w6481 & w6482) | (w6481 & w7788) | (w6482 & w7788);
assign w6484 = ~w6482 & w7789;
assign w6485 = ~w6483 & ~w6484;
assign w6486 = (~w6367 & ~w6369) | (~w6367 & w8881) | (~w6369 & w8881);
assign w6487 = pi22 & ~w2588;
assign w6488 = pi23 & w2390;
assign w6489 = (pi59 & w6487) | (pi59 & w8882) | (w6487 & w8882);
assign w6490 = ~w6487 & w8883;
assign w6491 = ~w6489 & ~w6490;
assign w6492 = pi18 & ~w3404;
assign w6493 = pi19 & w3186;
assign w6494 = (pi63 & w6492) | (pi63 & w7790) | (w6492 & w7790);
assign w6495 = ~w6492 & w7791;
assign w6496 = ~w6494 & ~w6495;
assign w6497 = pi20 & ~w2981;
assign w6498 = pi21 & w2932;
assign w6499 = (pi61 & w6497) | (pi61 & w7792) | (w6497 & w7792);
assign w6500 = ~w6497 & w7793;
assign w6501 = ~w6499 & ~w6500;
assign w6502 = w6496 & w6501;
assign w6503 = ~w6496 & ~w6501;
assign w6504 = ~w6502 & ~w6503;
assign w6505 = w6491 & w6504;
assign w6506 = ~w6491 & ~w6504;
assign w6507 = ~w6505 & ~w6506;
assign w6508 = ~w6486 & w6507;
assign w6509 = w6486 & ~w6507;
assign w6510 = ~w6508 & ~w6509;
assign w6511 = w6373 & w6510;
assign w6512 = ~w6373 & ~w6510;
assign w6513 = ~w6511 & ~w6512;
assign w6514 = ~w6432 & ~w6446;
assign w6515 = w6513 & w6514;
assign w6516 = ~w6513 & ~w6514;
assign w6517 = ~w6515 & ~w6516;
assign w6518 = w6395 & ~w6400;
assign w6519 = ~w6427 & ~w6518;
assign w6520 = pi30 & ~w1260;
assign w6521 = pi31 & ~w1131;
assign w6522 = ~w1130 & w6521;
assign w6523 = (pi51 & w6520) | (pi51 & w7948) | (w6520 & w7948);
assign w6524 = ~w6520 & w7949;
assign w6525 = ~w6523 & ~w6524;
assign w6526 = pi27 & w1695;
assign w6527 = pi26 & ~w1865;
assign w6528 = ~w1864 & w6527;
assign w6529 = ~w6526 & ~w6528;
assign w6530 = pi55 & ~w6529;
assign w6531 = ~pi55 & w6529;
assign w6532 = ~w6530 & ~w6531;
assign w6533 = pi29 & w1393;
assign w6534 = pi28 & ~w2050;
assign w6535 = ~w2049 & w6534;
assign w6536 = ~w6533 & ~w6535;
assign w6537 = pi53 & ~w6536;
assign w6538 = ~pi53 & w6536;
assign w6539 = ~w6537 & ~w6538;
assign w6540 = w6532 & w6539;
assign w6541 = ~w6532 & ~w6539;
assign w6542 = ~w6540 & ~w6541;
assign w6543 = w6525 & w6542;
assign w6544 = ~w6525 & ~w6542;
assign w6545 = ~w6543 & ~w6544;
assign w6546 = pi25 & w2032;
assign w6547 = pi24 & ~w2206;
assign w6548 = (pi57 & w6547) | (pi57 & w7950) | (w6547 & w7950);
assign w6549 = ~w6547 & w7951;
assign w6550 = ~w6548 & ~w6549;
assign w6551 = ~w6406 & ~w6422;
assign w6552 = (~w6550 & w6551) | (~w6550 & w7794) | (w6551 & w7794);
assign w6553 = ~w6551 & w7795;
assign w6554 = ~w6552 & ~w6553;
assign w6555 = ~w6545 & w6554;
assign w6556 = w6545 & ~w6554;
assign w6557 = ~w6555 & ~w6556;
assign w6558 = w6519 & w6557;
assign w6559 = ~w6519 & ~w6557;
assign w6560 = ~w6558 & ~w6559;
assign w6561 = ~w6438 & ~w6560;
assign w6562 = w6438 & w6560;
assign w6563 = ~w6561 & ~w6562;
assign w6564 = w6445 & w6563;
assign w6565 = ~w6445 & ~w6560;
assign w6566 = ~w6564 & ~w6565;
assign w6567 = w6517 & ~w6566;
assign w6568 = ~w6517 & w6566;
assign w6569 = ~w6567 & ~w6568;
assign w6570 = w6485 & ~w6569;
assign w6571 = ~w6485 & w6569;
assign w6572 = ~w6570 & ~w6571;
assign w6573 = w6480 & ~w6572;
assign w6574 = ~w6480 & w6572;
assign w6575 = ~w6573 & ~w6574;
assign w6576 = ~w6458 & ~w6575;
assign w6577 = w6458 & w6575;
assign w6578 = ~w6576 & ~w6577;
assign w6579 = ~w6476 & w7952;
assign w6580 = ~w6459 & ~w6575;
assign w6581 = w6459 & w6575;
assign w6582 = ~w6580 & ~w6581;
assign w6583 = (w6582 & w6476) | (w6582 & w7953) | (w6476 & w7953);
assign w6584 = ~w6579 & ~w6583;
assign w6585 = w6338 & w6460;
assign w6586 = w6214 & w6585;
assign w6587 = w6585 & w7954;
assign w6588 = w6462 & w6587;
assign w6589 = w6588 & w9087;
assign w6590 = w5648 & w6588;
assign w6591 = w5650 & w6590;
assign w6592 = (w6591 & w4814) | (w6591 & w7955) | (w4814 & w7955);
assign w6593 = ~w6589 & ~w6592;
assign w6594 = ~w6511 & ~w6515;
assign w6595 = ~w6517 & ~w6565;
assign w6596 = (w6594 & w6595) | (w6594 & w7796) | (w6595 & w7796);
assign w6597 = ~w6595 & w7797;
assign w6598 = ~w6596 & ~w6597;
assign w6599 = pi27 & ~w5754;
assign w6600 = (pi55 & w6599) | (pi55 & w7798) | (w6599 & w7798);
assign w6601 = ~w6599 & w7799;
assign w6602 = ~w6600 & ~w6601;
assign w6603 = pi29 & ~w1536;
assign w6604 = pi30 & w1393;
assign w6605 = (pi53 & w6603) | (pi53 & w7800) | (w6603 & w7800);
assign w6606 = ~w6603 & w7801;
assign w6607 = ~w6605 & ~w6606;
assign w6608 = w6602 & w6607;
assign w6609 = ~w6602 & ~w6607;
assign w6610 = ~w6608 & ~w6609;
assign w6611 = (pi51 & w1131) | (pi51 & w8885) | (w1131 & w8885);
assign w6612 = pi31 & ~pi51;
assign w6613 = ~w1130 & w6612;
assign w6614 = ~w6611 & ~w6613;
assign w6615 = ~w6610 & ~w6614;
assign w6616 = w6610 & w6614;
assign w6617 = ~w6615 & ~w6616;
assign w6618 = (~w6540 & ~w6542) | (~w6540 & w7802) | (~w6542 & w7802);
assign w6619 = pi25 & ~w2206;
assign w6620 = pi26 & w2032;
assign w6621 = (pi57 & w6619) | (pi57 & w8886) | (w6619 & w8886);
assign w6622 = ~w6619 & w8887;
assign w6623 = ~w6621 & ~w6622;
assign w6624 = w6618 & ~w6623;
assign w6625 = ~w6618 & w6623;
assign w6626 = ~w6624 & ~w6625;
assign w6627 = w6617 & ~w6626;
assign w6628 = ~w6617 & w6626;
assign w6629 = ~w6627 & ~w6628;
assign w6630 = ~w6552 & ~w6555;
assign w6631 = ~w6629 & w6630;
assign w6632 = w6629 & ~w6630;
assign w6633 = ~w6631 & ~w6632;
assign w6634 = (~w6502 & ~w6504) | (~w6502 & w8888) | (~w6504 & w8888);
assign w6635 = pi23 & ~w2588;
assign w6636 = pi24 & w2390;
assign w6637 = (pi59 & w6635) | (pi59 & w8889) | (w6635 & w8889);
assign w6638 = ~w6635 & w8890;
assign w6639 = ~w6637 & ~w6638;
assign w6640 = pi19 & ~w3404;
assign w6641 = (pi63 & w6640) | (pi63 & w7803) | (w6640 & w7803);
assign w6642 = ~w6640 & w7804;
assign w6643 = ~w6641 & ~w6642;
assign w6644 = pi21 & ~w2981;
assign w6645 = pi22 & w2932;
assign w6646 = (pi61 & w6644) | (pi61 & w7805) | (w6644 & w7805);
assign w6647 = ~w6644 & w7806;
assign w6648 = ~w6646 & ~w6647;
assign w6649 = w6643 & w6648;
assign w6650 = ~w6643 & ~w6648;
assign w6651 = ~w6649 & ~w6650;
assign w6652 = w6639 & w6651;
assign w6653 = ~w6639 & ~w6651;
assign w6654 = ~w6652 & ~w6653;
assign w6655 = ~w6634 & w6654;
assign w6656 = w6634 & ~w6654;
assign w6657 = ~w6655 & ~w6656;
assign w6658 = w6508 & w6657;
assign w6659 = ~w6508 & ~w6657;
assign w6660 = ~w6658 & ~w6659;
assign w6661 = w6438 & ~w6559;
assign w6662 = ~w6438 & ~w6558;
assign w6663 = ~w6661 & ~w6662;
assign w6664 = w6660 & ~w6663;
assign w6665 = ~w6660 & w6663;
assign w6666 = ~w6664 & ~w6665;
assign w6667 = w6633 & w6666;
assign w6668 = ~w6633 & ~w6666;
assign w6669 = ~w6667 & ~w6668;
assign w6670 = ~w6598 & ~w6669;
assign w6671 = w6598 & w6669;
assign w6672 = ~w6670 & ~w6671;
assign w6673 = ~w6484 & w6569;
assign w6674 = ~w6483 & ~w6673;
assign w6675 = w6672 & w6674;
assign w6676 = ~w6672 & ~w6674;
assign w6677 = ~w6675 & ~w6676;
assign w6678 = ~w6337 & ~w6459;
assign w6679 = ~w6458 & ~w6678;
assign w6680 = ~w6336 & w6460;
assign w6681 = w6460 & w7807;
assign w6682 = ~w6679 & ~w6681;
assign w6683 = w6215 & w6587;
assign w6684 = (~w6574 & w6682) | (~w6574 & w8006) | (w6682 & w8006);
assign w6685 = ~w6683 & w6684;
assign w6686 = w6677 & w6685;
assign w6687 = ~w6677 & ~w6685;
assign w6688 = ~w6686 & ~w6687;
assign w6689 = ~w6592 & w8041;
assign w6690 = (~w6677 & w6592) | (~w6677 & w8042) | (w6592 & w8042);
assign w6691 = ~w6689 & ~w6690;
assign w6692 = (~w6597 & ~w6598) | (~w6597 & w7956) | (~w6598 & w7956);
assign w6693 = w6563 & ~w6666;
assign w6694 = ~w6667 & ~w6693;
assign w6695 = pi28 & ~w5754;
assign w6696 = pi29 & w1695;
assign w6697 = (pi55 & w6695) | (pi55 & w8891) | (w6695 & w8891);
assign w6698 = ~w6695 & w8892;
assign w6699 = ~w6697 & ~w6698;
assign w6700 = pi30 & ~w1536;
assign w6701 = pi31 & ~w1392;
assign w6702 = ~w1391 & w6701;
assign w6703 = (pi53 & w6700) | (pi53 & w8893) | (w6700 & w8893);
assign w6704 = ~w6700 & w8894;
assign w6705 = ~w6703 & ~w6704;
assign w6706 = w6699 & w6705;
assign w6707 = ~w6699 & ~w6705;
assign w6708 = ~w6706 & ~w6707;
assign w6709 = (~w6608 & ~w6610) | (~w6608 & w7957) | (~w6610 & w7957);
assign w6710 = pi26 & ~w2206;
assign w6711 = pi27 & w2032;
assign w6712 = (pi57 & w6710) | (pi57 & w8895) | (w6710 & w8895);
assign w6713 = ~w6710 & w8896;
assign w6714 = ~w6712 & ~w6713;
assign w6715 = w6709 & ~w6714;
assign w6716 = ~w6709 & w6714;
assign w6717 = ~w6715 & ~w6716;
assign w6718 = w6708 & ~w6717;
assign w6719 = ~w6708 & w6717;
assign w6720 = ~w6718 & ~w6719;
assign w6721 = (~w6624 & ~w6626) | (~w6624 & w8897) | (~w6626 & w8897);
assign w6722 = w6720 & w6721;
assign w6723 = ~w6720 & ~w6721;
assign w6724 = ~w6722 & ~w6723;
assign w6725 = (~w6649 & ~w6651) | (~w6649 & w7958) | (~w6651 & w7958);
assign w6726 = pi24 & ~w2588;
assign w6727 = pi25 & w2390;
assign w6728 = (pi59 & w6726) | (pi59 & w8898) | (w6726 & w8898);
assign w6729 = ~w6726 & w8899;
assign w6730 = ~w6728 & ~w6729;
assign w6731 = pi20 & ~w3404;
assign w6732 = (pi63 & w6731) | (pi63 & w7808) | (w6731 & w7808);
assign w6733 = ~w6731 & w7809;
assign w6734 = ~w6732 & ~w6733;
assign w6735 = pi22 & ~w2981;
assign w6736 = (pi61 & w6735) | (pi61 & w7810) | (w6735 & w7810);
assign w6737 = ~w6735 & w7811;
assign w6738 = ~w6736 & ~w6737;
assign w6739 = w6734 & w6738;
assign w6740 = ~w6734 & ~w6738;
assign w6741 = ~w6739 & ~w6740;
assign w6742 = w6730 & w6741;
assign w6743 = ~w6730 & ~w6741;
assign w6744 = ~w6742 & ~w6743;
assign w6745 = w6725 & ~w6744;
assign w6746 = ~w6725 & w6744;
assign w6747 = ~w6745 & ~w6746;
assign w6748 = w6655 & w6747;
assign w6749 = ~w6655 & ~w6747;
assign w6750 = ~w6748 & ~w6749;
assign w6751 = w6631 & w6750;
assign w6752 = ~w6631 & ~w6750;
assign w6753 = ~w6751 & ~w6752;
assign w6754 = w6724 & w6753;
assign w6755 = ~w6724 & ~w6753;
assign w6756 = ~w6754 & ~w6755;
assign w6757 = ~w6559 & ~w6658;
assign w6758 = (~w6659 & w6562) | (~w6659 & w8900) | (w6562 & w8900);
assign w6759 = w6756 & w6758;
assign w6760 = ~w6756 & ~w6758;
assign w6761 = ~w6759 & ~w6760;
assign w6762 = ~w6694 & w6761;
assign w6763 = w6694 & ~w6761;
assign w6764 = ~w6762 & ~w6763;
assign w6765 = w6692 & ~w6764;
assign w6766 = ~w6692 & w6764;
assign w6767 = ~w6765 & ~w6766;
assign w6768 = w6685 & w8901;
assign w6769 = ~w6676 & w6767;
assign w6770 = w6676 & ~w6767;
assign w6771 = ~w6769 & ~w6770;
assign w6772 = (~w6771 & ~w6685) | (~w6771 & w8902) | (~w6685 & w8902);
assign w6773 = ~w6768 & ~w6772;
assign w6774 = ~w5949 & w6773;
assign w6775 = w6086 & w6587;
assign w6776 = w6685 & w8903;
assign w6777 = w6767 & w6776;
assign w6778 = w6771 & ~w6776;
assign w6779 = ~w6777 & ~w6778;
assign w6780 = w5949 & ~w6779;
assign w6781 = ~w6774 & ~w6780;
assign w6782 = w5946 & w6775;
assign w6783 = (w6782 & ~w5328) | (w6782 & w7959) | (~w5328 & w7959);
assign w6784 = w7738 & w8904;
assign w6785 = w6775 & w6784;
assign w6786 = ~w5333 & w6785;
assign w6787 = (~w7959 & w8905) | (~w7959 & w8906) | (w8905 & w8906);
assign w6788 = w6677 & w6767;
assign w6789 = w6575 & w6788;
assign w6790 = ~w5929 & ~w6080;
assign w6791 = w6586 & w7812;
assign w6792 = ~w5801 & w6791;
assign w6793 = ~w5937 & w6792;
assign w6794 = w5945 & w7813;
assign w6795 = w6791 & w6794;
assign w6796 = ~w6793 & ~w6795;
assign w6797 = pi29 & ~w5754;
assign w6798 = pi30 & w1695;
assign w6799 = (pi55 & w6797) | (pi55 & w8907) | (w6797 & w8907);
assign w6800 = ~w6797 & w8908;
assign w6801 = ~w6799 & ~w6800;
assign w6802 = (pi53 & w1392) | (pi53 & w8909) | (w1392 & w8909);
assign w6803 = pi31 & ~pi53;
assign w6804 = ~w1391 & w6803;
assign w6805 = ~w6802 & ~w6804;
assign w6806 = w6801 & w6805;
assign w6807 = ~w6801 & ~w6805;
assign w6808 = ~w6806 & ~w6807;
assign w6809 = pi27 & ~w2206;
assign w6810 = pi28 & w2032;
assign w6811 = (pi57 & w6809) | (pi57 & w8910) | (w6809 & w8910);
assign w6812 = ~w6809 & w8911;
assign w6813 = ~w6811 & ~w6812;
assign w6814 = w6707 & ~w6813;
assign w6815 = ~w6707 & w6813;
assign w6816 = ~w6814 & ~w6815;
assign w6817 = w6808 & w6816;
assign w6818 = ~w6808 & ~w6816;
assign w6819 = ~w6817 & ~w6818;
assign w6820 = (~w6716 & ~w6717) | (~w6716 & w8912) | (~w6717 & w8912);
assign w6821 = ~w6819 & w6820;
assign w6822 = w6819 & ~w6820;
assign w6823 = ~w6821 & ~w6822;
assign w6824 = (~w6739 & ~w6741) | (~w6739 & w8913) | (~w6741 & w8913);
assign w6825 = pi25 & ~w2588;
assign w6826 = pi26 & w2390;
assign w6827 = (pi59 & w6825) | (pi59 & w8914) | (w6825 & w8914);
assign w6828 = ~w6825 & w8915;
assign w6829 = ~w6827 & ~w6828;
assign w6830 = pi21 & ~w3404;
assign w6831 = pi22 & w3186;
assign w6832 = (pi63 & w6830) | (pi63 & w8043) | (w6830 & w8043);
assign w6833 = ~w6830 & w8044;
assign w6834 = ~w6832 & ~w6833;
assign w6835 = pi23 & ~w2981;
assign w6836 = pi24 & w2932;
assign w6837 = (pi61 & w6835) | (pi61 & w8045) | (w6835 & w8045);
assign w6838 = ~w6835 & w8046;
assign w6839 = ~w6837 & ~w6838;
assign w6840 = w6834 & w6839;
assign w6841 = ~w6834 & ~w6839;
assign w6842 = ~w6840 & ~w6841;
assign w6843 = w6829 & w6842;
assign w6844 = ~w6829 & ~w6842;
assign w6845 = ~w6843 & ~w6844;
assign w6846 = w6824 & ~w6845;
assign w6847 = ~w6824 & w6845;
assign w6848 = ~w6846 & ~w6847;
assign w6849 = w6746 & w6848;
assign w6850 = ~w6746 & ~w6848;
assign w6851 = ~w6849 & ~w6850;
assign w6852 = w6722 & w6851;
assign w6853 = ~w6722 & ~w6851;
assign w6854 = ~w6852 & ~w6853;
assign w6855 = ~w6823 & ~w6854;
assign w6856 = w6823 & w6854;
assign w6857 = ~w6855 & ~w6856;
assign w6858 = w6753 & w8916;
assign w6859 = (~w6748 & ~w6753) | (~w6748 & w8917) | (~w6753 & w8917);
assign w6860 = ~w6858 & ~w6859;
assign w6861 = ~w6751 & ~w6860;
assign w6862 = w6857 & ~w6861;
assign w6863 = ~w6857 & w6861;
assign w6864 = ~w6862 & ~w6863;
assign w6865 = (~w6759 & ~w6761) | (~w6759 & w8918) | (~w6761 & w8918);
assign w6866 = w6864 & ~w6865;
assign w6867 = ~w6864 & w6865;
assign w6868 = ~w6866 & ~w6867;
assign w6869 = ~w6675 & ~w6766;
assign w6870 = ~w6765 & ~w6869;
assign w6871 = (w6868 & w6869) | (w6868 & w8919) | (w6869 & w8919);
assign w6872 = ~w6869 & w8920;
assign w6873 = ~w6871 & ~w6872;
assign w6874 = w6796 & w8921;
assign w6875 = w6788 & ~w6873;
assign w6876 = ~w6788 & w6873;
assign w6877 = ~w6875 & ~w6876;
assign w6878 = (~w6877 & ~w6796) | (~w6877 & w8922) | (~w6796 & w8922);
assign w6879 = ~w6874 & ~w6878;
assign w6880 = w6787 & ~w6879;
assign w6881 = (~w6877 & w6783) | (~w6877 & w8047) | (w6783 & w8047);
assign w6882 = ~w6880 & ~w6881;
assign w6883 = ~w6788 & ~w6870;
assign w6884 = ~w6574 & ~w6870;
assign w6885 = (w6884 & w6682) | (w6884 & w7960) | (w6682 & w7960);
assign w6886 = ~w6683 & w6885;
assign w6887 = ~w6883 & ~w6886;
assign w6888 = ~w6792 & ~w6887;
assign w6889 = w5320 & w5940;
assign w6890 = w4998 & w6889;
assign w6891 = ~w6888 & w6890;
assign w6892 = ~w4237 & w6891;
assign w6893 = w4993 & w6889;
assign w6894 = w5942 & ~w6887;
assign w6895 = (~w6888 & ~w6894) | (~w6888 & w7961) | (~w6894 & w7961);
assign w6896 = (~w6858 & w6861) | (~w6858 & w8923) | (w6861 & w8923);
assign w6897 = (~w6815 & ~w6816) | (~w6815 & w8924) | (~w6816 & w8924);
assign w6898 = pi30 & ~w5754;
assign w6899 = pi31 & ~w1694;
assign w6900 = ~w1693 & w6899;
assign w6901 = (pi55 & w6898) | (pi55 & w8925) | (w6898 & w8925);
assign w6902 = ~w6898 & w8926;
assign w6903 = ~w6901 & ~w6902;
assign w6904 = pi28 & ~w2206;
assign w6905 = pi29 & w2032;
assign w6906 = (pi57 & w6904) | (pi57 & w8927) | (w6904 & w8927);
assign w6907 = ~w6904 & w8928;
assign w6908 = ~w6906 & ~w6907;
assign w6909 = w6806 & w6908;
assign w6910 = ~w6806 & ~w6908;
assign w6911 = ~w6909 & ~w6910;
assign w6912 = ~w6903 & w6911;
assign w6913 = w6903 & ~w6911;
assign w6914 = ~w6912 & ~w6913;
assign w6915 = w6897 & ~w6914;
assign w6916 = ~w6897 & w6914;
assign w6917 = ~w6915 & ~w6916;
assign w6918 = (~w6840 & ~w6842) | (~w6840 & w8929) | (~w6842 & w8929);
assign w6919 = pi26 & ~w2588;
assign w6920 = pi27 & w2390;
assign w6921 = (pi59 & w6919) | (pi59 & w8930) | (w6919 & w8930);
assign w6922 = ~w6919 & w8931;
assign w6923 = ~w6921 & ~w6922;
assign w6924 = pi22 & ~w3404;
assign w6925 = pi23 & w3186;
assign w6926 = (pi63 & w6924) | (pi63 & w8932) | (w6924 & w8932);
assign w6927 = ~w6924 & w8933;
assign w6928 = ~w6926 & ~w6927;
assign w6929 = pi24 & ~w2981;
assign w6930 = pi25 & w2932;
assign w6931 = (pi61 & w6929) | (pi61 & w8934) | (w6929 & w8934);
assign w6932 = ~w6929 & w8935;
assign w6933 = ~w6931 & ~w6932;
assign w6934 = w6928 & w6933;
assign w6935 = ~w6928 & ~w6933;
assign w6936 = ~w6934 & ~w6935;
assign w6937 = w6923 & w6936;
assign w6938 = ~w6923 & ~w6936;
assign w6939 = ~w6937 & ~w6938;
assign w6940 = w6918 & ~w6939;
assign w6941 = ~w6918 & w6939;
assign w6942 = ~w6940 & ~w6941;
assign w6943 = w6847 & w6942;
assign w6944 = ~w6847 & ~w6942;
assign w6945 = ~w6943 & ~w6944;
assign w6946 = w6822 & w6945;
assign w6947 = ~w6822 & ~w6945;
assign w6948 = ~w6946 & ~w6947;
assign w6949 = w6917 & w6948;
assign w6950 = ~w6917 & ~w6948;
assign w6951 = ~w6949 & ~w6950;
assign w6952 = w6854 & w8936;
assign w6953 = (~w6849 & ~w6854) | (~w6849 & w8937) | (~w6854 & w8937);
assign w6954 = ~w6952 & ~w6953;
assign w6955 = ~w6852 & ~w6954;
assign w6956 = w6951 & ~w6955;
assign w6957 = ~w6951 & w6955;
assign w6958 = ~w6956 & ~w6957;
assign w6959 = ~w6896 & w6958;
assign w6960 = w6896 & ~w6958;
assign w6961 = ~w6959 & ~w6960;
assign w6962 = ~w6867 & w6961;
assign w6963 = w6867 & ~w6961;
assign w6964 = w6866 & w6961;
assign w6965 = ~w6866 & ~w6961;
assign w6966 = ~w6892 & w8048;
assign w6967 = ~w6963 & ~w6964;
assign w6968 = (~w6892 & w8959) | (~w6892 & w8960) | (w8959 & w8960);
assign w6969 = ~w6966 & w6968;
assign w6970 = (~w6909 & ~w6911) | (~w6909 & w8938) | (~w6911 & w8938);
assign w6971 = pi29 & ~w2206;
assign w6972 = pi30 & w2032;
assign w6973 = (pi57 & w6971) | (pi57 & w8939) | (w6971 & w8939);
assign w6974 = ~w6971 & w8940;
assign w6975 = ~w6973 & ~w6974;
assign w6976 = w6903 & w6975;
assign w6977 = ~w6903 & ~w6975;
assign w6978 = ~w6976 & ~w6977;
assign w6979 = (pi55 & w1694) | (pi55 & w8941) | (w1694 & w8941);
assign w6980 = pi31 & ~pi55;
assign w6981 = ~w1693 & w6980;
assign w6982 = ~w6979 & ~w6981;
assign w6983 = ~w6978 & ~w6982;
assign w6984 = w6978 & w6982;
assign w6985 = ~w6983 & ~w6984;
assign w6986 = ~w6970 & w6985;
assign w6987 = w6970 & ~w6985;
assign w6988 = ~w6986 & ~w6987;
assign w6989 = (~w6934 & ~w6936) | (~w6934 & w8942) | (~w6936 & w8942);
assign w6990 = pi27 & ~w2588;
assign w6991 = pi28 & w2390;
assign w6992 = (pi59 & w6990) | (pi59 & w8943) | (w6990 & w8943);
assign w6993 = ~w6990 & w8944;
assign w6994 = ~w6992 & ~w6993;
assign w6995 = pi23 & ~w3404;
assign w6996 = pi24 & w3186;
assign w6997 = (pi63 & w6995) | (pi63 & w8945) | (w6995 & w8945);
assign w6998 = ~w6995 & w8946;
assign w6999 = ~w6997 & ~w6998;
assign w7000 = pi25 & ~w2981;
assign w7001 = pi26 & w2932;
assign w7002 = (pi61 & w7000) | (pi61 & w8947) | (w7000 & w8947);
assign w7003 = ~w7000 & w8948;
assign w7004 = ~w7002 & ~w7003;
assign w7005 = w6999 & w7004;
assign w7006 = ~w6999 & ~w7004;
assign w7007 = ~w7005 & ~w7006;
assign w7008 = w6994 & w7007;
assign w7009 = ~w6994 & ~w7007;
assign w7010 = ~w7008 & ~w7009;
assign w7011 = w6989 & ~w7010;
assign w7012 = ~w6989 & w7010;
assign w7013 = ~w7011 & ~w7012;
assign w7014 = w6941 & w7013;
assign w7015 = ~w6941 & ~w7013;
assign w7016 = ~w7014 & ~w7015;
assign w7017 = w6916 & w7016;
assign w7018 = ~w6916 & ~w7016;
assign w7019 = ~w7017 & ~w7018;
assign w7020 = w6988 & w7019;
assign w7021 = ~w6988 & ~w7019;
assign w7022 = ~w7020 & ~w7021;
assign w7023 = w6948 & w8949;
assign w7024 = (~w6943 & ~w6948) | (~w6943 & w8961) | (~w6948 & w8961);
assign w7025 = ~w7023 & ~w7024;
assign w7026 = ~w6946 & ~w7025;
assign w7027 = w7022 & ~w7026;
assign w7028 = ~w7022 & w7026;
assign w7029 = ~w7027 & ~w7028;
assign w7030 = ~w6952 & ~w6956;
assign w7031 = ~w7029 & w7030;
assign w7032 = w7029 & ~w7030;
assign w7033 = ~w7031 & ~w7032;
assign w7034 = ~w6883 & ~w6884;
assign w7035 = w6459 & w6789;
assign w7036 = ~w7034 & ~w7035;
assign w7037 = ~w6867 & ~w6960;
assign w7038 = (~w6959 & ~w6961) | (~w6959 & w8962) | (~w6961 & w8962);
assign w7039 = (w7038 & w7036) | (w7038 & w8049) | (w7036 & w8049);
assign w7040 = w6868 & w6961;
assign w7041 = w6680 & w6789;
assign w7042 = w7040 & w7041;
assign w7043 = w7039 & ~w7042;
assign w7044 = (w6469 & w7963) | (w6469 & w7964) | (w7963 & w7964);
assign w7045 = (~w6469 & w7965) | (~w6469 & w7966) | (w7965 & w7966);
assign w7046 = ~w7044 & ~w7045;
assign w7047 = ~w7023 & ~w7027;
assign w7048 = ~w6976 & ~w6984;
assign w7049 = pi30 & ~w2206;
assign w7050 = pi31 & w2032;
assign w7051 = ~w7049 & ~w7050;
assign w7052 = pi57 & ~w7051;
assign w7053 = ~pi57 & w7051;
assign w7054 = ~w7052 & ~w7053;
assign w7055 = w7048 & w7054;
assign w7056 = ~w7048 & ~w7054;
assign w7057 = ~w7055 & ~w7056;
assign w7058 = (~w7005 & ~w7007) | (~w7005 & w7814) | (~w7007 & w7814);
assign w7059 = pi28 & ~w2588;
assign w7060 = pi29 & w2390;
assign w7061 = ~w7059 & ~w7060;
assign w7062 = pi59 & ~w7061;
assign w7063 = ~pi59 & w7061;
assign w7064 = ~w7062 & ~w7063;
assign w7065 = pi24 & ~w3404;
assign w7066 = (pi63 & w7065) | (pi63 & w7815) | (w7065 & w7815);
assign w7067 = ~w7065 & w7816;
assign w7068 = ~w7066 & ~w7067;
assign w7069 = pi26 & ~w2981;
assign w7070 = pi27 & w2932;
assign w7071 = (pi61 & w7069) | (pi61 & w7817) | (w7069 & w7817);
assign w7072 = ~w7069 & w7818;
assign w7073 = ~w7071 & ~w7072;
assign w7074 = w7068 & w7073;
assign w7075 = ~w7068 & ~w7073;
assign w7076 = ~w7074 & ~w7075;
assign w7077 = w7064 & w7076;
assign w7078 = ~w7064 & ~w7076;
assign w7079 = ~w7077 & ~w7078;
assign w7080 = w7058 & ~w7079;
assign w7081 = ~w7058 & w7079;
assign w7082 = ~w7080 & ~w7081;
assign w7083 = w7012 & w7082;
assign w7084 = ~w7012 & ~w7082;
assign w7085 = ~w7083 & ~w7084;
assign w7086 = w6986 & w7085;
assign w7087 = ~w6986 & ~w7085;
assign w7088 = ~w7086 & ~w7087;
assign w7089 = w7057 & w7088;
assign w7090 = ~w7057 & ~w7088;
assign w7091 = ~w7089 & ~w7090;
assign w7092 = w7019 & w7819;
assign w7093 = (~w7014 & ~w7019) | (~w7014 & w7820) | (~w7019 & w7820);
assign w7094 = ~w7092 & ~w7093;
assign w7095 = ~w7017 & ~w7094;
assign w7096 = w7091 & ~w7095;
assign w7097 = ~w7091 & w7095;
assign w7098 = ~w7096 & ~w7097;
assign w7099 = ~w7047 & w7098;
assign w7100 = w7047 & ~w7098;
assign w7101 = ~w7099 & ~w7100;
assign w7102 = ~w7031 & w7101;
assign w7103 = w7031 & ~w7101;
assign w7104 = ~w7102 & ~w7103;
assign w7105 = (~w6469 & w7967) | (~w6469 & w7968) | (w7967 & w7968);
assign w7106 = ~w7033 & w7104;
assign w7107 = w7033 & w7101;
assign w7108 = ~w7106 & ~w7107;
assign w7109 = (w6469 & w7969) | (w6469 & w7970) | (w7969 & w7970);
assign w7110 = ~w7105 & ~w7109;
assign w7111 = pi31 & ~w2031;
assign w7112 = pi57 & ~w7111;
assign w7113 = pi31 & ~pi57;
assign w7114 = ~w2030 & w7113;
assign w7115 = ~w7112 & ~w7114;
assign w7116 = w7054 & w7115;
assign w7117 = ~w7054 & ~w7115;
assign w7118 = ~w7116 & ~w7117;
assign w7119 = (~w7074 & ~w7076) | (~w7074 & w8963) | (~w7076 & w8963);
assign w7120 = pi29 & ~w2588;
assign w7121 = pi30 & w2390;
assign w7122 = ~w7120 & ~w7121;
assign w7123 = pi59 & ~w7122;
assign w7124 = ~pi59 & w7122;
assign w7125 = ~w7123 & ~w7124;
assign w7126 = pi25 & ~w3404;
assign w7127 = (pi63 & w7126) | (pi63 & w7821) | (w7126 & w7821);
assign w7128 = ~w7126 & w7822;
assign w7129 = ~w7127 & ~w7128;
assign w7130 = pi27 & ~w2981;
assign w7131 = pi28 & w2932;
assign w7132 = (pi61 & w7130) | (pi61 & w7823) | (w7130 & w7823);
assign w7133 = ~w7130 & w7824;
assign w7134 = ~w7132 & ~w7133;
assign w7135 = w7129 & w7134;
assign w7136 = ~w7129 & ~w7134;
assign w7137 = ~w7135 & ~w7136;
assign w7138 = w7125 & w7137;
assign w7139 = ~w7125 & ~w7137;
assign w7140 = ~w7138 & ~w7139;
assign w7141 = w7119 & ~w7140;
assign w7142 = ~w7119 & w7140;
assign w7143 = ~w7141 & ~w7142;
assign w7144 = w7081 & w7143;
assign w7145 = ~w7081 & ~w7143;
assign w7146 = ~w7144 & ~w7145;
assign w7147 = w7056 & w7146;
assign w7148 = ~w7056 & ~w7146;
assign w7149 = ~w7147 & ~w7148;
assign w7150 = ~w7118 & ~w7149;
assign w7151 = w7118 & w7149;
assign w7152 = ~w7150 & ~w7151;
assign w7153 = w7088 & w8964;
assign w7154 = (~w7083 & ~w7088) | (~w7083 & w8965) | (~w7088 & w8965);
assign w7155 = ~w7153 & ~w7154;
assign w7156 = ~w7086 & ~w7155;
assign w7157 = w7152 & ~w7156;
assign w7158 = ~w7152 & w7156;
assign w7159 = ~w7157 & ~w7158;
assign w7160 = ~w7092 & ~w7096;
assign w7161 = ~w7159 & w7160;
assign w7162 = w7159 & ~w7160;
assign w7163 = ~w7161 & ~w7162;
assign w7164 = w7040 & w7107;
assign w7165 = w6789 & w7164;
assign w7166 = w6585 & w7165;
assign w7167 = w5650 & w8966;
assign w7168 = (w7167 & w4814) | (w7167 & w8050) | (w4814 & w8050);
assign w7169 = ~w6585 & ~w6679;
assign w7170 = ~w5656 & w7825;
assign w7171 = ~w6471 & w8051;
assign w7172 = ~w6473 & w7171;
assign w7173 = w7165 & ~w7169;
assign w7174 = (w7173 & w7170) | (w7173 & w8052) | (w7170 & w8052);
assign w7175 = w7034 & w7164;
assign w7176 = ~w7032 & ~w7099;
assign w7177 = ~w7100 & ~w7176;
assign w7178 = ~w7038 & w7102;
assign w7179 = ~w7177 & ~w7178;
assign w7180 = ~w7175 & w7179;
assign w7181 = (w7163 & w7168) | (w7163 & w7826) | (w7168 & w7826);
assign w7182 = ~w7168 & w7827;
assign w7183 = ~w7181 & ~w7182;
assign w7184 = w7163 & w7179;
assign w7185 = (w7184 & w6886) | (w7184 & w8967) | (w6886 & w8967);
assign w7186 = ~w7165 & w7185;
assign w7187 = ~w7153 & ~w7157;
assign w7188 = w7149 & w8968;
assign w7189 = (~w7144 & ~w7149) | (~w7144 & w8969) | (~w7149 & w8969);
assign w7190 = ~w7188 & ~w7189;
assign w7191 = ~w7147 & ~w7190;
assign w7192 = ~w7135 & ~w7138;
assign w7193 = pi30 & ~w2588;
assign w7194 = pi31 & w2390;
assign w7195 = ~w7193 & ~w7194;
assign w7196 = pi59 & ~w7195;
assign w7197 = ~pi59 & w7195;
assign w7198 = ~w7196 & ~w7197;
assign w7199 = pi26 & ~w3404;
assign w7200 = pi27 & w3186;
assign w7201 = ~w7199 & ~w7200;
assign w7202 = pi63 & ~w7201;
assign w7203 = ~pi63 & w7201;
assign w7204 = ~w7202 & ~w7203;
assign w7205 = pi28 & ~w2981;
assign w7206 = pi29 & w2932;
assign w7207 = ~w7205 & ~w7206;
assign w7208 = pi61 & ~w7207;
assign w7209 = ~pi61 & w7207;
assign w7210 = ~w7208 & ~w7209;
assign w7211 = w7204 & w7210;
assign w7212 = ~w7204 & ~w7210;
assign w7213 = ~w7211 & ~w7212;
assign w7214 = w7198 & w7213;
assign w7215 = ~w7198 & ~w7213;
assign w7216 = ~w7214 & ~w7215;
assign w7217 = w7192 & ~w7216;
assign w7218 = ~w7192 & w7216;
assign w7219 = ~w7217 & ~w7218;
assign w7220 = w7142 & w7219;
assign w7221 = ~w7142 & ~w7219;
assign w7222 = ~w7220 & ~w7221;
assign w7223 = w7116 & ~w7222;
assign w7224 = ~w7116 & w7222;
assign w7225 = ~w7223 & ~w7224;
assign w7226 = w7191 & ~w7225;
assign w7227 = ~w7191 & w7225;
assign w7228 = ~w7226 & ~w7227;
assign w7229 = ~w7187 & w7228;
assign w7230 = w7187 & ~w7228;
assign w7231 = ~w7229 & ~w7230;
assign w7232 = ~w7161 & w7231;
assign w7233 = w7161 & ~w7231;
assign w7234 = ~w7232 & ~w7233;
assign w7235 = ~w7186 & ~w7234;
assign w7236 = w7186 & w7234;
assign w7237 = ~w7235 & ~w7236;
assign w7238 = ~w6593 & w7237;
assign w7239 = ~w7185 & ~w7234;
assign w7240 = w7185 & w7234;
assign w7241 = ~w7239 & ~w7240;
assign w7242 = ~w6592 & w7829;
assign w7243 = ~w7238 & ~w7242;
assign w7244 = ~w7188 & ~w7227;
assign w7245 = ~w7116 & w7221;
assign w7246 = w7116 & w7220;
assign w7247 = ~w7245 & ~w7246;
assign w7248 = ~w7211 & ~w7214;
assign w7249 = pi27 & ~w3404;
assign w7250 = pi28 & w3186;
assign w7251 = ~w7249 & ~w7250;
assign w7252 = pi63 & ~w7251;
assign w7253 = ~pi63 & w7251;
assign w7254 = ~w7252 & ~w7253;
assign w7255 = pi29 & ~w2981;
assign w7256 = pi30 & w2932;
assign w7257 = ~w7255 & ~w7256;
assign w7258 = pi61 & ~w7257;
assign w7259 = ~pi61 & w7257;
assign w7260 = ~w7258 & ~w7259;
assign w7261 = w7254 & w7260;
assign w7262 = ~w7254 & ~w7260;
assign w7263 = ~w7261 & ~w7262;
assign w7264 = pi31 & ~w2389;
assign w7265 = pi59 & ~w7264;
assign w7266 = pi31 & ~pi59;
assign w7267 = ~w2388 & w7266;
assign w7268 = ~w7265 & ~w7267;
assign w7269 = ~w7263 & ~w7268;
assign w7270 = w7263 & w7268;
assign w7271 = ~w7269 & ~w7270;
assign w7272 = w7248 & ~w7271;
assign w7273 = ~w7248 & w7271;
assign w7274 = ~w7272 & ~w7273;
assign w7275 = ~w7218 & ~w7274;
assign w7276 = w7218 & w7274;
assign w7277 = ~w7275 & ~w7276;
assign w7278 = w7247 & ~w7277;
assign w7279 = ~w7247 & w7277;
assign w7280 = ~w7278 & ~w7279;
assign w7281 = ~w7244 & ~w7280;
assign w7282 = w7244 & w7280;
assign w7283 = ~w7281 & ~w7282;
assign w7284 = ~w7161 & ~w7230;
assign w7285 = ~w7229 & ~w7284;
assign w7286 = w6588 & w7165;
assign w7287 = w6784 & w7286;
assign w7288 = ~w7162 & ~w7229;
assign w7289 = w7179 & w7288;
assign w7290 = (w7289 & w5333) | (w7289 & w8970) | (w5333 & w8970);
assign w7291 = w7167 & ~w7285;
assign w7292 = (w7291 & ~w5328) | (w7291 & w8053) | (~w5328 & w8053);
assign w7293 = (w7283 & w7292) | (w7283 & w7971) | (w7292 & w7971);
assign w7294 = ~w7292 & w7972;
assign w7295 = ~w7293 & ~w7294;
assign w7296 = w7283 & ~w7285;
assign w7297 = ~w7289 & w7296;
assign w7298 = w7164 & w7296;
assign w7299 = ~w7297 & w7298;
assign w7300 = ~w7245 & ~w7278;
assign w7301 = ~w7261 & ~w7270;
assign w7302 = pi28 & ~w3404;
assign w7303 = pi29 & w3186;
assign w7304 = ~w7302 & ~w7303;
assign w7305 = pi63 & ~w7304;
assign w7306 = ~pi63 & w7304;
assign w7307 = ~w7305 & ~w7306;
assign w7308 = pi30 & ~w2981;
assign w7309 = pi31 & w2932;
assign w7310 = ~w7308 & ~w7309;
assign w7311 = pi61 & ~w7310;
assign w7312 = ~pi61 & w7310;
assign w7313 = ~w7311 & ~w7312;
assign w7314 = w7307 & w7313;
assign w7315 = ~w7307 & ~w7313;
assign w7316 = ~w7314 & ~w7315;
assign w7317 = ~w7301 & ~w7316;
assign w7318 = w7301 & w7316;
assign w7319 = ~w7317 & ~w7318;
assign w7320 = ~w7273 & ~w7276;
assign w7321 = w7319 & ~w7320;
assign w7322 = ~w7319 & w7320;
assign w7323 = ~w7321 & ~w7322;
assign w7324 = w7300 & w7323;
assign w7325 = ~w7300 & ~w7323;
assign w7326 = ~w7324 & ~w7325;
assign w7327 = ~w7281 & ~w7297;
assign w7328 = w7326 & ~w7327;
assign w7329 = ~w7326 & w7327;
assign w7330 = ~w7328 & ~w7329;
assign w7331 = (w7830 & w6892) | (w7830 & w8953) | (w6892 & w8953);
assign w7332 = (~w6892 & w8954) | (~w6892 & w8955) | (w8954 & w8955);
assign w7333 = ~w7331 & ~w7332;
assign w7334 = w7276 & w7319;
assign w7335 = pi29 & ~w3404;
assign w7336 = pi30 & w3186;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = pi63 & ~w7337;
assign w7339 = ~pi63 & w7337;
assign w7340 = ~w7338 & ~w7339;
assign w7341 = pi31 & ~w2931;
assign w7342 = pi61 & ~w7341;
assign w7343 = pi31 & ~pi61;
assign w7344 = ~w2930 & w7343;
assign w7345 = ~w7342 & ~w7344;
assign w7346 = w7340 & w7345;
assign w7347 = ~w7340 & ~w7345;
assign w7348 = ~w7346 & ~w7347;
assign w7349 = w7315 & ~w7348;
assign w7350 = ~w7315 & w7348;
assign w7351 = ~w7349 & ~w7350;
assign w7352 = w7273 & w7319;
assign w7353 = ~w7317 & ~w7352;
assign w7354 = w7351 & ~w7353;
assign w7355 = ~w7351 & w7353;
assign w7356 = ~w7354 & ~w7355;
assign w7357 = w7334 & w7356;
assign w7358 = ~w7334 & ~w7356;
assign w7359 = ~w7357 & ~w7358;
assign w7360 = ~w7282 & w7326;
assign w7361 = w7162 & ~w7230;
assign w7362 = ~w7229 & ~w7281;
assign w7363 = ~w7361 & w7362;
assign w7364 = w7284 & w7360;
assign w7365 = w7363 & w7364;
assign w7366 = w7107 & w7365;
assign w7367 = w7359 & w7366;
assign w7368 = w7360 & ~w7363;
assign w7369 = ~w7324 & ~w7368;
assign w7370 = w7177 & w7365;
assign w7371 = w7369 & ~w7370;
assign w7372 = w7359 & ~w7371;
assign w7373 = ~w7359 & w7371;
assign w7374 = ~w7372 & ~w7373;
assign w7375 = ~w7366 & ~w7374;
assign w7376 = ~w7367 & ~w7375;
assign w7377 = (~w6469 & w7973) | (~w6469 & w7974) | (w7973 & w7974);
assign w7378 = (w6469 & w7975) | (w6469 & w7976) | (w7975 & w7976);
assign w7379 = ~w7377 & ~w7378;
assign w7380 = w6462 & w7832;
assign w7381 = w7041 & w8971;
assign w7382 = (w7381 & ~w6472) | (w7381 & w7833) | (~w6472 & w7833);
assign w7383 = ~w7357 & w7371;
assign w7384 = (w7383 & w7039) | (w7383 & w7834) | (w7039 & w7834);
assign w7385 = ~w7382 & w7384;
assign w7386 = ~w7358 & w7365;
assign w7387 = w5939 & w7386;
assign w7388 = w7286 & w7387;
assign w7389 = ~w7382 & w8956;
assign w7390 = (w7389 & w5651) | (w7389 & w7977) | (w5651 & w7977);
assign w7391 = w7351 & w7352;
assign w7392 = w7317 & w7351;
assign w7393 = pi30 & ~w3404;
assign w7394 = pi31 & w3186;
assign w7395 = ~w7393 & ~w7394;
assign w7396 = pi63 & ~w7395;
assign w7397 = ~pi63 & w7395;
assign w7398 = ~w7396 & ~w7397;
assign w7399 = ~w7346 & ~w7350;
assign w7400 = w7398 & ~w7399;
assign w7401 = ~w7398 & w7399;
assign w7402 = ~w7400 & ~w7401;
assign w7403 = w7392 & ~w7402;
assign w7404 = ~w7392 & w7402;
assign w7405 = ~w7403 & ~w7404;
assign w7406 = w7391 & w7405;
assign w7407 = ~w7391 & ~w7405;
assign w7408 = ~w7406 & ~w7407;
assign w7409 = ~w7385 & w7978;
assign w7410 = (w7408 & w7385) | (w7408 & w7979) | (w7385 & w7979);
assign w7411 = ~w7409 & ~w7410;
assign w7412 = w7390 & w7411;
assign w7413 = ~w7390 & ~w7411;
assign w7414 = ~w7412 & ~w7413;
assign w7415 = (~w7174 & w4821) | (~w7174 & w7835) | (w4821 & w7835);
assign w7416 = ~w7346 & ~w7398;
assign w7417 = pi31 & ~w3185;
assign w7418 = pi63 & ~w7417;
assign w7419 = pi31 & ~pi63;
assign w7420 = ~w3184 & w7419;
assign w7421 = ~w7418 & ~w7420;
assign w7422 = ~w7416 & w7421;
assign w7423 = w7416 & ~w7421;
assign w7424 = ~w7422 & ~w7423;
assign w7425 = w7350 & ~w7398;
assign w7426 = ~w7403 & ~w7425;
assign w7427 = w7424 & ~w7426;
assign w7428 = ~w7424 & w7426;
assign w7429 = ~w7427 & ~w7428;
assign w7430 = (~w7358 & w7368) | (~w7358 & w7980) | (w7368 & w7980);
assign w7431 = ~w7357 & ~w7406;
assign w7432 = ~w7430 & w7431;
assign w7433 = ~w7407 & ~w7432;
assign w7434 = w7180 & ~w7433;
assign w7435 = w7359 & w7408;
assign w7436 = w7365 & w7435;
assign w7437 = w7434 & w7436;
assign w7438 = w7429 & w7437;
assign w7439 = ~w7433 & ~w7436;
assign w7440 = w7429 & w7439;
assign w7441 = ~w7429 & ~w7439;
assign w7442 = ~w7440 & ~w7441;
assign w7443 = ~w7437 & ~w7442;
assign w7444 = ~w7438 & ~w7443;
assign w7445 = w7415 & ~w7444;
assign w7446 = ~w7442 & ~w7415;
assign w7447 = ~w7445 & ~w7446;
assign w7448 = w7423 & w7426;
assign w7449 = ~w7439 & ~w7448;
assign w7450 = ~w7422 & ~w7427;
assign w7451 = ~w7449 & w7450;
assign w7452 = w7434 & w7450;
assign w7453 = (w4821 & w8054) | (w4821 & w8055) | (w8054 & w8055);
assign w7454 = ~w7451 & ~w7453;
assign w7455 = w50 & pi35;
assign w7456 = ~w50 & ~pi35;
assign w7457 = ~pi02 & pi35;
assign w7458 = ~pi00 & pi37;
assign w7459 = ~w96 & w120;
assign w7460 = w96 & ~w120;
assign w7461 = ~pi03 & pi35;
assign w7462 = ~pi01 & pi37;
assign w7463 = w169 & pi39;
assign w7464 = ~w169 & ~pi39;
assign w7465 = ~pi04 & pi35;
assign w7466 = ~pi02 & pi37;
assign w7467 = w220 & pi39;
assign w7468 = ~w220 & ~pi39;
assign w7469 = ~pi05 & pi35;
assign w7470 = ~pi03 & pi37;
assign w7471 = ~w229 & w274;
assign w7472 = w229 & ~w274;
assign w7473 = ~pi35 & pi06;
assign w7474 = ~w283 & ~w289;
assign w7475 = w283 & w289;
assign w7476 = w306 & pi41;
assign w7477 = ~w306 & ~pi41;
assign w7478 = w311 & pi39;
assign w7479 = ~w311 & ~pi39;
assign w7480 = w321 & ~w347;
assign w7481 = ~w321 & w347;
assign w7482 = ~pi01 & pi41;
assign w7483 = w331 & w418;
assign w7484 = ~w331 & ~w418;
assign w7485 = ~pi02 & pi41;
assign w7486 = ~pi00 & pi43;
assign w7487 = w402 & ~w394;
assign w7488 = ~pi06 & pi37;
assign w7489 = ~pi08 & pi35;
assign w7490 = w352 & w481;
assign w7491 = w351 & w345;
assign w7492 = ~w351 & w494;
assign w7493 = ~w477 & ~w451;
assign w7494 = w474 & ~w466;
assign w7495 = ~pi01 & pi43;
assign w7496 = ~pi03 & pi41;
assign w7497 = ~pi07 & pi37;
assign w7498 = ~pi09 & pi35;
assign w7499 = ~w599 & w598;
assign w7500 = w54 & ~pi37;
assign w7501 = w8 & w7836;
assign w7502 = (~pi35 & ~w8) | (~pi35 & w7837) | (~w8 & w7837);
assign w7503 = ~pi02 & pi43;
assign w7504 = ~pi04 & pi41;
assign w7505 = w580 & ~w572;
assign w7506 = (~w692 & ~w622) | (~w692 & w7838) | (~w622 & w7838);
assign w7507 = w622 & w7839;
assign w7508 = ~w647 & ~w672;
assign w7509 = w217 & w7840;
assign w7510 = (~pi41 & ~w217) | (~pi41 & w7841) | (~w217 & w7841);
assign w7511 = w748 & pi35;
assign w7512 = ~w748 & ~pi35;
assign w7513 = w523 & w7981;
assign w7514 = (~pi45 & ~w523) | (~pi45 & w7982) | (~w523 & w7982);
assign w7515 = w856 & pi47;
assign w7516 = (~pi47 & ~w700) | (~pi47 & w7983) | (~w700 & w7983);
assign w7517 = w903 & pi45;
assign w7518 = ~w903 & ~pi45;
assign w7519 = ~w843 & ~w818;
assign w7520 = w840 & ~w832;
assign w7521 = w937 & pi39;
assign w7522 = ~w937 & ~pi39;
assign w7523 = w933 & w1009;
assign w7524 = ~w933 & ~w1009;
assign w7525 = w523 & w8972;
assign w7526 = (~pi45 & ~w523) | (~pi45 & w8973) | (~w523 & w8973);
assign w7527 = w982 & ~w974;
assign w7528 = w119 & w8974;
assign w7529 = (~pi39 & ~w119) | (~pi39 & w8975) | (~w119 & w8975);
assign w7530 = w523 & w9076;
assign w7531 = (~pi45 & ~w523) | (~pi45 & w8976) | (~w523 & w8976);
assign w7532 = w1097 & ~w1089;
assign w7533 = w119 & w8977;
assign w7534 = (~pi39 & ~w119) | (~pi39 & w8978) | (~w119 & w8978);
assign w7535 = ~w1137 & ~w1135;
assign w7536 = w1282 & pi45;
assign w7537 = ~w1282 & ~pi45;
assign w7538 = w1226 & ~w1218;
assign w7539 = w1314 & pi39;
assign w7540 = ~w1314 & ~pi39;
assign w7541 = ~w1268 & ~w1266;
assign w7542 = w523 & w8979;
assign w7543 = (~pi45 & ~w523) | (~pi45 & w8980) | (~w523 & w8980);
assign w7544 = w1359 & ~w1351;
assign w7545 = w119 & w8981;
assign w7546 = (~pi39 & ~w119) | (~pi39 & w8982) | (~w119 & w8982);
assign w7547 = ~w1414 & w7984;
assign w7548 = (~w1529 & w1414) | (~w1529 & w7985) | (w1414 & w7985);
assign w7549 = w1538 & pi53;
assign w7550 = ~w1538 & ~pi53;
assign w7551 = w1543 & pi51;
assign w7552 = ~w1543 & ~pi51;
assign w7553 = w1507 & ~w1453;
assign w7554 = w1501 & ~w1493;
assign w7555 = ~w1559 & w1557;
assign w7556 = ~w1559 & ~w1556;
assign w7557 = w1624 & ~w1616;
assign w7558 = ~w1533 & ~w1532;
assign w7559 = ~w1731 & w1851;
assign w7560 = w1731 & ~w1851;
assign w7561 = w1712 & ~w1705;
assign w7562 = w1857 & pi51;
assign w7563 = ~w1857 & ~pi51;
assign w7564 = ~w1718 & ~w1716;
assign w7565 = w1794 & ~w1786;
assign w7566 = w2042 & pi51;
assign w7567 = ~w2042 & ~pi51;
assign w7568 = w2092 & pi45;
assign w7569 = ~w2092 & ~pi45;
assign w7570 = w1961 & ~w1953;
assign w7571 = w2128 & pi39;
assign w7572 = ~w2128 & ~pi39;
assign w7573 = w2163 & w2169;
assign w7574 = ~w2163 & ~w2169;
assign w7575 = w2078 & w8983;
assign w7576 = (w2197 & ~w2078) | (w2197 & w8984) | (~w2078 & w8984);
assign w7577 = w2203 & pi57;
assign w7578 = ~w2203 & ~pi57;
assign w7579 = w2218 & pi51;
assign w7580 = ~w2218 & ~pi51;
assign w7581 = ~w2126 & w2175;
assign w7582 = w2266 & pi45;
assign w7583 = ~w2266 & ~pi45;
assign w7584 = w2301 & pi39;
assign w7585 = ~w2301 & ~pi39;
assign w7586 = w8 & w8985;
assign w7587 = (~pi35 & ~w8) | (~pi35 & w8986) | (~w8 & w8986);
assign w7588 = w56 & w9077;
assign w7589 = (~pi37 & ~w56) | (~pi37 & w8987) | (~w56 & w8987);
assign w7590 = ~w2023 & ~w2021;
assign w7591 = ~w2235 & w2411;
assign w7592 = ~pi03 & pi55;
assign w7593 = ~pi11 & pi47;
assign w7594 = ~pi17 & pi41;
assign w7595 = ~pi21 & pi37;
assign w7596 = ~pi23 & pi35;
assign w7597 = w2360 & ~w2363;
assign w7598 = w2253 & w2393;
assign w7599 = w2395 & ~w2393;
assign w7600 = ~w2433 & w2612;
assign w7601 = ~pi04 & pi55;
assign w7602 = ~pi10 & pi49;
assign w7603 = w2547 & ~w2539;
assign w7604 = ~pi16 & pi43;
assign w7605 = ~w2453 & w2594;
assign w7606 = ~w2596 & ~w2594;
assign w7607 = ~w2631 & w2786;
assign w7608 = ~pi05 & pi55;
assign w7609 = ~pi11 & pi49;
assign w7610 = w2715 & ~w2707;
assign w7611 = (w2974 & ~w2952) | (w2974 & w7842) | (~w2952 & w7842);
assign w7612 = w2952 & w7843;
assign w7613 = w2926 & ~w2826;
assign w7614 = ~w2805 & w3017;
assign w7615 = w2889 & ~w2881;
assign w7616 = ~w2761 & ~w2962;
assign w7617 = ~w2963 & ~w3171;
assign w7618 = ~w3036 & w3233;
assign w7619 = w3120 & ~w3112;
assign w7620 = w3220 & w7844;
assign w7621 = (w3391 & ~w3220) | (w3391 & w7845) | (~w3220 & w7845);
assign w7622 = ~w3252 & w3446;
assign w7623 = w3336 & ~w3328;
assign w7624 = ~w3606 & ~w3604;
assign w7625 = ~w3433 & w7846;
assign w7626 = (~w3621 & w3433) | (~w3621 & w7847) | (w3433 & w7847);
assign w7627 = ~w3465 & w3672;
assign w7628 = w3534 & ~w3547;
assign w7629 = w3659 & w7848;
assign w7630 = (~w3830 & ~w3659) | (~w3830 & w7849) | (~w3659 & w7849);
assign w7631 = w3842 & pi63;
assign w7632 = ~w3842 & ~pi63;
assign w7633 = w3847 & pi61;
assign w7634 = ~w3847 & ~pi61;
assign w7635 = ~w3691 & w3882;
assign w7636 = w3691 & ~w3882;
assign w7637 = w3963 & pi35;
assign w7638 = ~w3963 & ~pi35;
assign w7639 = w3968 & pi37;
assign w7640 = ~w3968 & ~pi37;
assign w7641 = w3755 & ~w3774;
assign w7642 = w3977 & pi39;
assign w7643 = ~w3977 & ~pi39;
assign w7644 = w3868 & w7986;
assign w7645 = (w4027 & ~w3868) | (w4027 & w7987) | (~w3868 & w7987);
assign w7646 = w4040 & pi63;
assign w7647 = ~w4040 & ~pi63;
assign w7648 = w4045 & pi61;
assign w7649 = ~w4045 & ~pi61;
assign w7650 = w3918 & w4065;
assign w7651 = ~w3900 & w4074;
assign w7652 = w3900 & ~w4074;
assign w7653 = w3884 & ~w3885;
assign w7654 = w3975 & ~w3974;
assign w7655 = ~pi31 & pi35;
assign w7656 = ~pi37 & ~w4174;
assign w7657 = w2371 & w2013;
assign w7658 = w4260 & pi63;
assign w7659 = ~w4260 & ~pi63;
assign w7660 = w4265 & pi61;
assign w7661 = ~w4265 & ~pi61;
assign w7662 = w4117 & ~w4285;
assign w7663 = ~w4092 & w4294;
assign w7664 = w4092 & ~w4294;
assign w7665 = ~w4181 & ~w4180;
assign w7666 = ~pi37 & ~pi30;
assign w7667 = w4347 & pi39;
assign w7668 = ~w4347 & ~pi39;
assign w7669 = w4385 & pi45;
assign w7670 = ~w4385 & ~pi45;
assign w7671 = w4156 & ~w4209;
assign w7672 = w4408 & ~w4382;
assign w7673 = ~w4350 & ~w4344;
assign w7674 = ~w4288 & w4614;
assign w7675 = w4472 & w4466;
assign w7676 = ~w4497 & w4651;
assign w7677 = w4497 & ~w4651;
assign w7678 = w4656 & pi51;
assign w7679 = ~w4656 & ~pi51;
assign w7680 = ~w4689 & ~w4576;
assign w7681 = w4517 & ~w4599;
assign w7682 = w4637 & ~w4804;
assign w7683 = ~w4637 & w4804;
assign w7684 = ~w3607 & w4813;
assign w7685 = w4653 & ~w4654;
assign w7686 = ~w4673 & w4842;
assign w7687 = ~w4721 & ~w4719;
assign w7688 = w4625 & ~w4809;
assign w7689 = ~w4992 & ~w4808;
assign w7690 = w3607 & w4995;
assign w7691 = ~w4874 & ~w4836;
assign w7692 = ~w4902 & ~w4900;
assign w7693 = ~w4860 & w5118;
assign w7694 = ~w5159 & ~w5009;
assign w7695 = w5047 & w7850;
assign w7696 = (~w5170 & ~w5047) | (~w5170 & w7851) | (~w5047 & w7851);
assign w7697 = w5150 & ~w5112;
assign w7698 = w5153 & ~w5106;
assign w7699 = ~w5136 & w5220;
assign w7700 = ~w5324 & ~w5327;
assign w7701 = (~w4989 & ~w4810) | (~w4989 & w7852) | (~w4810 & w7852);
assign w7702 = ~w5239 & w5349;
assign w7703 = w5206 & ~w5200;
assign w7704 = ~w5206 & ~w5485;
assign w7705 = w5478 & w5472;
assign w7706 = w5382 & ~w5343;
assign w7707 = ~w5368 & w5561;
assign w7708 = w5567 & pi51;
assign w7709 = ~w5567 & ~pi51;
assign w7710 = ~w5398 & ~w5411;
assign w7711 = w5642 & w5511;
assign w7712 = w5547 & w7988;
assign w7713 = (~w5665 & ~w5547) | (~w5665 & w7989) | (~w5547 & w7989);
assign w7714 = ~w5594 & ~w5554;
assign w7715 = w909 & w7853;
assign w7716 = (~pi49 & ~w909) | (~pi49 & w7854) | (~w909 & w7854);
assign w7717 = w5720 & pi47;
assign w7718 = (~pi47 & ~w700) | (~pi47 & w7855) | (~w700 & w7855);
assign w7719 = w5741 & pi57;
assign w7720 = ~w5741 & ~pi57;
assign w7721 = w5752 & pi55;
assign w7722 = ~w5752 & ~pi55;
assign w7723 = w5701 & ~w5810;
assign w7724 = ~w5701 & w5810;
assign w7725 = w5787 & ~w5783;
assign w7726 = ~w5773 & w5855;
assign w7727 = w5773 & ~w5855;
assign w7728 = w5860 & pi51;
assign w7729 = ~w5860 & ~pi51;
assign w7730 = w909 & w7856;
assign w7731 = (~pi49 & ~w909) | (~pi49 & w7857) | (~w909 & w7857);
assign w7732 = w700 & w7990;
assign w7733 = (~pi47 & ~w700) | (~pi47 & w7858) | (~w700 & w7858);
assign w7734 = ~w5738 & w5918;
assign w7735 = w5738 & ~w5918;
assign w7736 = w5668 & ~w5667;
assign w7737 = w5646 & ~w5800;
assign w7738 = w5649 & w5165;
assign w7739 = w5924 & ~w5812;
assign w7740 = w5738 & ~w5846;
assign w7741 = w5973 & pi63;
assign w7742 = ~w5973 & ~pi63;
assign w7743 = w5978 & pi61;
assign w7744 = ~w5978 & ~pi61;
assign w7745 = w6000 & pi57;
assign w7746 = ~w6000 & ~pi57;
assign w7747 = w6011 & pi51;
assign w7748 = ~w6011 & ~pi51;
assign w7749 = w5858 & ~w5857;
assign w7750 = w6107 & pi57;
assign w7751 = ~w6107 & ~pi57;
assign w7752 = w6118 & pi55;
assign w7753 = ~w6118 & ~pi55;
assign w7754 = w6150 & pi49;
assign w7755 = ~w6150 & ~pi49;
assign w7756 = w6180 & pi63;
assign w7757 = ~w6180 & ~pi63;
assign w7758 = w6185 & pi61;
assign w7759 = ~w6185 & ~pi61;
assign w7760 = ~w6039 & w5910;
assign w7761 = w6081 & ~w6080;
assign w7762 = ~w6171 & w6223;
assign w7763 = w6171 & ~w6223;
assign w7764 = w6239 & pi63;
assign w7765 = ~w6239 & ~pi63;
assign w7766 = w6244 & pi61;
assign w7767 = ~w6244 & ~pi61;
assign w7768 = ~w6137 & w6269;
assign w7769 = w6137 & ~w6269;
assign w7770 = w6274 & pi51;
assign w7771 = ~w6274 & ~pi51;
assign w7772 = w6321 & w6231;
assign w7773 = w6358 & pi63;
assign w7774 = ~w6358 & ~pi63;
assign w7775 = w6363 & pi61;
assign w7776 = ~w6363 & ~pi61;
assign w7777 = ~w6302 & ~w6162;
assign w7778 = w6391 & pi57;
assign w7779 = ~w6391 & ~pi57;
assign w7780 = w6402 & pi51;
assign w7781 = ~w6402 & ~pi51;
assign w7782 = w6272 & ~w6271;
assign w7783 = w6430 & ~w6311;
assign w7784 = ~w6311 & ~w6440;
assign w7785 = ~w6227 & ~w6225;
assign w7786 = w6461 & w5800;
assign w7787 = ~w6468 & w6475;
assign w7788 = ~w6386 & w7859;
assign w7789 = (~w6481 & w6386) | (~w6481 & w7860) | (w6386 & w7860);
assign w7790 = w6493 & pi63;
assign w7791 = ~w6493 & ~pi63;
assign w7792 = w6498 & pi61;
assign w7793 = ~w6498 & ~pi61;
assign w7794 = w6421 & ~w6550;
assign w7795 = ~w6421 & w6550;
assign w7796 = w6564 & w6594;
assign w7797 = ~w6564 & ~w6594;
assign w7798 = w1695 & w7861;
assign w7799 = (~pi55 & ~w1695) | (~pi55 & w7862) | (~w1695 & w7862);
assign w7800 = w6604 & pi53;
assign w7801 = (~pi53 & ~w1393) | (~pi53 & w7863) | (~w1393 & w7863);
assign w7802 = ~w6525 & ~w6540;
assign w7803 = w3186 & w7864;
assign w7804 = (~pi63 & ~w3186) | (~pi63 & w7865) | (~w3186 & w7865);
assign w7805 = w6645 & pi61;
assign w7806 = (~pi61 & ~w2932) | (~pi61 & w7866) | (~w2932 & w7866);
assign w7807 = ~w6336 & w6212;
assign w7808 = w3186 & w7867;
assign w7809 = (~pi63 & ~w3186) | (~pi63 & w7868) | (~w3186 & w7868);
assign w7810 = w2932 & w7991;
assign w7811 = (~pi61 & ~w2932) | (~pi61 & w7869) | (~w2932 & w7869);
assign w7812 = w6790 & w6789;
assign w7813 = w5497 & w8988;
assign w7814 = ~w6994 & ~w7005;
assign w7815 = w3186 & w7992;
assign w7816 = (~pi63 & ~w3186) | (~pi63 & w7993) | (~w3186 & w7993);
assign w7817 = w7070 & pi61;
assign w7818 = (~pi61 & ~w2932) | (~pi61 & w7994) | (~w2932 & w7994);
assign w7819 = w6988 & w7014;
assign w7820 = ~w6988 & ~w7014;
assign w7821 = w3186 & w7995;
assign w7822 = (~pi63 & ~w3186) | (~pi63 & w7996) | (~w3186 & w7996);
assign w7823 = w7131 & pi61;
assign w7824 = (~pi61 & ~w2932) | (~pi61 & w7997) | (~w2932 & w7997);
assign w7825 = w5932 & w6463;
assign w7826 = (w7163 & w7174) | (w7163 & w7998) | (w7174 & w7998);
assign w7827 = ~w7174 & w7999;
assign w7828 = ~w6883 & w7164;
assign w7829 = ~w6589 & w7241;
assign w7830 = w7299 & w7330;
assign w7831 = ~w7299 & ~w7330;
assign w7832 = ~w5800 & w5647;
assign w7833 = w7380 & w7381;
assign w7834 = w7371 & w8000;
assign w7835 = ~w7167 & ~w7174;
assign w7836 = pi11 & pi35;
assign w7837 = ~pi11 & ~pi35;
assign w7838 = w620 & ~w692;
assign w7839 = ~w620 & w692;
assign w7840 = pi06 & pi41;
assign w7841 = ~pi06 & ~pi41;
assign w7842 = ~w2950 & w2974;
assign w7843 = w2950 & ~w2974;
assign w7844 = w3218 & ~w3391;
assign w7845 = ~w3218 & w3391;
assign w7846 = ~w3431 & w3621;
assign w7847 = w3431 & ~w3621;
assign w7848 = ~w3657 & w3830;
assign w7849 = w3657 & ~w3830;
assign w7850 = ~w5045 & w5170;
assign w7851 = w5045 & ~w5170;
assign w7852 = ~w4020 & ~w4989;
assign w7853 = pi27 & pi49;
assign w7854 = ~pi27 & ~pi49;
assign w7855 = ~pi29 & ~pi47;
assign w7856 = pi28 & pi49;
assign w7857 = ~pi28 & ~pi49;
assign w7858 = ~pi30 & ~pi47;
assign w7859 = ~w6385 & w6481;
assign w7860 = w6385 & ~w6481;
assign w7861 = pi28 & pi55;
assign w7862 = ~pi28 & ~pi55;
assign w7863 = ~pi30 & ~pi53;
assign w7864 = pi20 & pi63;
assign w7865 = ~pi20 & ~pi63;
assign w7866 = ~pi22 & ~pi61;
assign w7867 = pi21 & pi63;
assign w7868 = ~pi21 & ~pi63;
assign w7869 = ~pi23 & ~pi61;
assign w7870 = ~w7039 & ~w7043;
assign w7871 = ~w496 & ~w493;
assign w7872 = ~w528 & ~w527;
assign w7873 = w523 & w8001;
assign w7874 = (~pi45 & ~w523) | (~pi45 & w8002) | (~w523 & w8002);
assign w7875 = w644 & ~w636;
assign w7876 = ~w711 & ~w709;
assign w7877 = w873 & w896;
assign w7878 = ~w873 & ~w896;
assign w7879 = w900 & w895;
assign w7880 = ~w900 & w1111;
assign w7881 = ~w1120 & ~w1117;
assign w7882 = ~w1246 & w1520;
assign w7883 = w1559 & w1556;
assign w7884 = w1845 & w1520;
assign w7885 = ~w1839 & ~w2006;
assign w7886 = ~w2011 & ~w2377;
assign w7887 = w2374 & ~w2382;
assign w7888 = ~w3003 & ~w3001;
assign w7889 = ~w2382 & ~w3600;
assign w7890 = w3385 & ~w3597;
assign w7891 = w3615 & ~w4234;
assign w7892 = w4239 & w4224;
assign w7893 = w4291 & pi57;
assign w7894 = ~w4291 & ~pi57;
assign w7895 = w3607 & w4629;
assign w7896 = ~w4815 & ~w4819;
assign w7897 = (~w4827 & ~w4798) | (~w4827 & w8989) | (~w4798 & w8989);
assign w7898 = w4798 & w8990;
assign w7899 = w4224 & w4810;
assign w7900 = ~w4999 & ~w4994;
assign w7901 = ~w4831 & ~w4829;
assign w7902 = w5022 & pi63;
assign w7903 = ~w5022 & ~pi63;
assign w7904 = w5027 & pi61;
assign w7905 = ~w5027 & ~pi61;
assign w7906 = w4860 & ~w5118;
assign w7907 = w5182 & pi63;
assign w7908 = ~w5182 & ~pi63;
assign w7909 = w5187 & pi61;
assign w7910 = ~w5187 & ~pi61;
assign w7911 = w5120 & ~w5121;
assign w7912 = w4810 & w4021;
assign w7913 = w4224 & w4022;
assign w7914 = ~w3611 & w5324;
assign w7915 = w4224 & w3823;
assign w7916 = (w5319 & w8003) | (w5319 & w9093) | (w8003 & w9093);
assign w7917 = ~w5202 & ~w5200;
assign w7918 = w4815 & w5650;
assign w7919 = w5163 & ~w5317;
assign w7920 = ~w5653 & ~w5496;
assign w7921 = ~w5660 & w5648;
assign w7922 = w5678 & pi63;
assign w7923 = ~w5678 & ~pi63;
assign w7924 = w5683 & pi61;
assign w7925 = ~w5683 & ~pi61;
assign w7926 = w5627 & ~w5431;
assign w7927 = w5824 & pi63;
assign w7928 = ~w5824 & ~pi63;
assign w7929 = w5829 & pi61;
assign w7930 = ~w5829 & ~pi61;
assign w7931 = w5852 & pi57;
assign w7932 = ~w5852 & ~pi57;
assign w7933 = ~w5712 & ~w5724;
assign w7934 = ~w5944 & ~w5948;
assign w7935 = ~w5844 & ~w5842;
assign w7936 = ~w5738 & w5962;
assign w7937 = ~w5906 & ~w5900;
assign w7938 = w6076 & w5958;
assign w7939 = ~w6071 & w6095;
assign w7940 = w6071 & ~w6095;
assign w7941 = ~w6092 & w6218;
assign w7942 = w6091 & w6339;
assign w7943 = ~w6218 & w8004;
assign w7944 = (~w6338 & w6218) | (~w6338 & w8005) | (w6218 & w8005);
assign w7945 = w6461 & ~w5800;
assign w7946 = w6336 & w6460;
assign w7947 = ~w6336 & ~w6460;
assign w7948 = w6522 & pi51;
assign w7949 = ~w6522 & ~pi51;
assign w7950 = w6546 & pi57;
assign w7951 = ~w6546 & ~pi57;
assign w7952 = ~w6336 & ~w6578;
assign w7953 = w6336 & w6582;
assign w7954 = w6214 & w6575;
assign w7955 = ~w4820 & w6591;
assign w7956 = ~w6669 & ~w6597;
assign w7957 = ~w6614 & ~w6608;
assign w7958 = ~w6639 & ~w6649;
assign w7959 = w7914 & w8991;
assign w7960 = ~w6870 & w8006;
assign w7961 = w6893 & ~w6888;
assign w7962 = (w7961 & w8957) | (w7961 & w8958) | (w8957 & w8958);
assign w7963 = w7033 & w7043;
assign w7964 = (w6475 & w7963) | (w6475 & w8007) | (w7963 & w8007);
assign w7965 = ~w7033 & ~w7043;
assign w7966 = ~w7033 & w9094;
assign w7967 = ~w7104 & ~w7043;
assign w7968 = ~w7104 & w9094;
assign w7969 = w7108 & w7043;
assign w7970 = (w6475 & w7969) | (w6475 & w8008) | (w7969 & w8008);
assign w7971 = (~w7290 & w7296) | (~w7290 & w8057) | (w7296 & w8057);
assign w7972 = (w7290 & w8011) | (w7290 & w8012) | (w8011 & w8012);
assign w7973 = ~w7376 & ~w7043;
assign w7974 = ~w7376 & w9094;
assign w7975 = ~w7374 & w7043;
assign w7976 = (w6475 & w7975) | (w6475 & w8013) | (w7975 & w8013);
assign w7977 = ~w5660 & w7389;
assign w7978 = ~w7358 & ~w7408;
assign w7979 = w7358 & w7408;
assign w7980 = w7324 & ~w7358;
assign w7981 = pi03 & pi45;
assign w7982 = ~pi03 & ~pi45;
assign w7983 = ~pi01 & ~pi47;
assign w7984 = ~w1412 & w1529;
assign w7985 = w1412 & ~w1529;
assign w7986 = w3866 & ~w4027;
assign w7987 = ~w3866 & w4027;
assign w7988 = ~w5546 & w5665;
assign w7989 = w5546 & ~w5665;
assign w7990 = pi30 & pi47;
assign w7991 = pi23 & pi61;
assign w7992 = pi25 & pi63;
assign w7993 = ~pi25 & ~pi63;
assign w7994 = ~pi27 & ~pi61;
assign w7995 = pi26 & pi63;
assign w7996 = ~pi26 & ~pi63;
assign w7997 = ~pi28 & ~pi61;
assign w7998 = ~w7180 & w7163;
assign w7999 = w7180 & ~w7163;
assign w8000 = ~w7357 & ~w7366;
assign w8001 = pi02 & pi45;
assign w8002 = ~pi02 & ~pi45;
assign w8003 = w5331 & w5319;
assign w8004 = w6339 & w6338;
assign w8005 = ~w6339 & ~w6338;
assign w8006 = ~w6574 & w6573;
assign w8007 = w7033 & ~w7870;
assign w8008 = w7108 & ~w7870;
assign w8009 = ~w7285 & w7164;
assign w8010 = ~w6886 & w8992;
assign w8011 = ~w7283 & w7285;
assign w8012 = (w6796 & w8993) | (w6796 & w8994) | (w8993 & w8994);
assign w8013 = ~w7374 & ~w7870;
assign w8014 = ~w720 & ~w731;
assign w8015 = ~w701 & ~w863;
assign w8016 = w847 & ~w865;
assign w8017 = ~w1106 & ~w1012;
assign w8018 = ~w2371 & ~w2572;
assign w8019 = ~w3175 & ~w3173;
assign w8020 = ~w4022 & ~w3823;
assign w8021 = ~w4434 & ~w4224;
assign w8022 = ~w4434 & ~w7892;
assign w8023 = ~w4631 & ~w4431;
assign w8024 = ~w4989 & ~w4994;
assign w8025 = ~w4989 & w7900;
assign w8026 = w5335 & ~w5319;
assign w8027 = w5501 & ~w5319;
assign w8028 = w5501 & ~w7916;
assign w8029 = w4810 & w5649;
assign w8030 = w5660 & ~w5648;
assign w8031 = w5801 & ~w5947;
assign w8032 = w5946 & w6086;
assign w8033 = ~w6214 & ~w6212;
assign w8034 = w7943 & w6338;
assign w8035 = (w6338 & w7943) | (w6338 & w6340) | (w7943 & w6340);
assign w8036 = ~w6340 & w7944;
assign w8037 = ~w3607 & w6466;
assign w8038 = w5650 & w8995;
assign w8039 = ~w6337 & w6339;
assign w8040 = ~w6470 & w6474;
assign w8041 = ~w6589 & ~w6688;
assign w8042 = w6589 & ~w6677;
assign w8043 = w6831 & pi63;
assign w8044 = ~w6831 & ~pi63;
assign w8045 = w6836 & pi61;
assign w8046 = ~w6836 & ~pi61;
assign w8047 = w6786 & ~w6877;
assign w8048 = w6965 & ~w6895;
assign w8049 = ~w7037 & w7038;
assign w8050 = ~w4820 & w7167;
assign w8051 = w6339 & ~w6679;
assign w8052 = ~w7172 & w7173;
assign w8053 = w5325 & w7291;
assign w8054 = w7452 & ~w7174;
assign w8055 = w7452 & w7835;
assign w8056 = ~w6091 & w6093;
assign w8057 = w7283 & w9095;
assign w8058 = w6216 & ~w6093;
assign w8059 = w6216 & w9088;
assign w8060 = w17 & w11;
assign w8061 = w27 & pi35;
assign w8062 = ~w27 & ~pi35;
assign w8063 = ~pi00 & pi35;
assign w8064 = ~w9 & ~w40;
assign w8065 = ~w22 & ~w42;
assign w8066 = pi00 & ~pi37;
assign w8067 = ~w36 & pi37;
assign w8068 = w36 & ~pi37;
assign w8069 = w68 & ~w60;
assign w8070 = ~pi35 & pi02;
assign w8071 = ~w83 & ~w84;
assign w8072 = ~w89 & ~w91;
assign w8073 = ~w74 & ~w72;
assign w8074 = ~pi35 & pi03;
assign w8075 = ~w126 & ~w127;
assign w8076 = ~pi37 & pi01;
assign w8077 = ~w132 & ~w133;
assign w8078 = ~w107 & ~w151;
assign w8079 = ~pi00 & pi39;
assign w8080 = ~w96 & w158;
assign w8081 = ~pi35 & pi04;
assign w8082 = ~w180 & ~w181;
assign w8083 = ~pi37 & pi02;
assign w8084 = ~w186 & ~w187;
assign w8085 = ~w153 & ~w208;
assign w8086 = ~pi35 & pi05;
assign w8087 = ~w233 & ~w234;
assign w8088 = ~pi37 & pi03;
assign w8089 = ~w239 & ~w240;
assign w8090 = ~pi00 & pi41;
assign w8091 = ~w218 & ~w273;
assign w8092 = ~pi06 & pi35;
assign w8093 = ~w280 & ~w281;
assign w8094 = ~pi04 & pi37;
assign w8095 = pi05 & pi37;
assign w8096 = w295 & ~w297;
assign w8097 = w298 & ~w291;
assign w8098 = pi00 & ~pi43;
assign w8099 = ~pi41 & pi01;
assign w8100 = ~w360 & ~w361;
assign w8101 = w369 & pi39;
assign w8102 = ~w369 & ~pi39;
assign w8103 = ~pi05 & ~pi37;
assign w8104 = w426 & pi39;
assign w8105 = ~w426 & ~pi39;
assign w8106 = ~pi41 & pi02;
assign w8107 = ~w431 & ~w432;
assign w8108 = pi41 & pi00;
assign w8109 = ~w437 & ~w440;
assign w8110 = ~pi37 & pi06;
assign w8111 = ~w455 & ~w456;
assign w8112 = ~pi35 & pi08;
assign w8113 = ~w461 & ~w462;
assign w8114 = w372 & ~w366;
assign w8115 = w375 & ~w366;
assign w8116 = ~w375 & ~w481;
assign w8117 = w375 & w486;
assign w8118 = ~w415 & ~w500;
assign w8119 = w487 & ~w481;
assign w8120 = w480 & ~w519;
assign w8121 = ~w429 & ~w444;
assign w8122 = w535 & pi39;
assign w8123 = ~w535 & ~pi39;
assign w8124 = pi41 & pi01;
assign w8125 = ~w540 & ~w541;
assign w8126 = ~pi41 & pi03;
assign w8127 = ~w546 & ~w547;
assign w8128 = ~pi37 & pi07;
assign w8129 = ~w561 & ~w562;
assign w8130 = ~pi35 & pi09;
assign w8131 = ~w567 & ~w568;
assign w8132 = w599 & ~w598;
assign w8133 = w538 & ~w551;
assign w8134 = pi00 & pi45;
assign w8135 = w523 & w9089;
assign w8136 = ~w614 & ~w609;
assign w8137 = w557 & w620;
assign w8138 = ~w557 & ~w620;
assign w8139 = w649 & pi39;
assign w8140 = ~w649 & ~pi39;
assign w8141 = pi41 & pi02;
assign w8142 = ~w654 & ~w655;
assign w8143 = ~pi41 & pi04;
assign w8144 = ~w660 & ~w661;
assign w8145 = w590 & w683;
assign w8146 = ~w590 & ~w683;
assign w8147 = w597 & w686;
assign w8148 = ~w597 & ~w686;
assign w8149 = ~pi00 & pi45;
assign w8150 = ~w614 & w690;
assign w8151 = ~w652 & ~w665;
assign w8152 = w717 & pi39;
assign w8153 = ~w717 & ~pi39;
assign w8154 = ~pi03 & pi43;
assign w8155 = ~w727 & ~w726;
assign w8156 = ~w680 & ~w606;
assign w8157 = ~w684 & ~w686;
assign w8158 = ~w684 & ~w8147;
assign w8159 = w776 & ~w8157;
assign w8160 = w776 & ~w8158;
assign w8161 = ~w714 & w709;
assign w8162 = w714 & w781;
assign w8163 = w785 & pi39;
assign w8164 = ~w785 & ~pi39;
assign w8165 = ~pi10 & pi37;
assign w8166 = ~w822 & ~w821;
assign w8167 = ~pi12 & pi35;
assign w8168 = ~w828 & ~w827;
assign w8169 = ~pi00 & pi47;
assign w8170 = ~w774 & w885;
assign w8171 = w774 & ~w885;
assign w8172 = w776 & ~w685;
assign w8173 = ~w783 & ~w780;
assign w8174 = ~w788 & ~w809;
assign w8175 = ~pi00 & pi49;
assign w8176 = pi00 & ~pi49;
assign w8177 = ~pi01 & pi47;
assign w8178 = ~w915 & ~w914;
assign w8179 = ~pi07 & pi41;
assign w8180 = ~w943 & ~w942;
assign w8181 = ~pi05 & pi43;
assign w8182 = ~w949 & ~w948;
assign w8183 = ~pi13 & pi35;
assign w8184 = ~w964 & ~w963;
assign w8185 = ~pi11 & pi37;
assign w8186 = ~w970 & ~w969;
assign w8187 = ~w891 & ~w1002;
assign w8188 = ~pi02 & pi47;
assign w8189 = ~w1027 & ~w1026;
assign w8190 = ~w1033 & ~w1032;
assign w8191 = ~pi08 & pi41;
assign w8192 = ~w1058 & ~w1057;
assign w8193 = ~pi06 & pi43;
assign w8194 = ~w1064 & ~w1063;
assign w8195 = ~pi12 & pi37;
assign w8196 = ~w1079 & ~w1078;
assign w8197 = ~pi14 & pi35;
assign w8198 = ~w1085 & ~w1084;
assign w8199 = w997 & ~w884;
assign w8200 = w890 & ~w1121;
assign w8201 = ~w1042 & ~w1018;
assign w8202 = w1049 & ~w1137;
assign w8203 = ~w1049 & w1137;
assign w8204 = ~pi03 & pi47;
assign w8205 = ~w1156 & ~w1155;
assign w8206 = ~pi01 & pi49;
assign w8207 = ~w1162 & ~w1161;
assign w8208 = ~pi09 & pi41;
assign w8209 = ~w1187 & ~w1186;
assign w8210 = ~pi07 & pi43;
assign w8211 = ~w1193 & ~w1192;
assign w8212 = ~pi15 & pi35;
assign w8213 = ~w1208 & ~w1207;
assign w8214 = ~pi13 & pi37;
assign w8215 = ~w1214 & ~w1213;
assign w8216 = ~w1109 & ~w1110;
assign w8217 = w890 & w1246;
assign w8218 = ~w1140 & w1135;
assign w8219 = ~w1171 & ~w1147;
assign w8220 = pi00 & pi51;
assign w8221 = w1132 & w9090;
assign w8222 = ~w1262 & ~w1257;
assign w8223 = w1178 & ~w1268;
assign w8224 = ~w1178 & w1268;
assign w8225 = ~pi04 & pi47;
assign w8226 = ~w1288 & ~w1287;
assign w8227 = ~pi02 & pi49;
assign w8228 = ~w1294 & ~w1293;
assign w8229 = ~pi10 & pi41;
assign w8230 = ~w1320 & ~w1319;
assign w8231 = ~pi08 & pi43;
assign w8232 = ~w1326 & ~w1325;
assign w8233 = ~pi14 & pi37;
assign w8234 = ~w1341 & ~w1340;
assign w8235 = ~pi16 & pi35;
assign w8236 = ~w1347 & ~w1346;
assign w8237 = ~w1380 & ~w1379;
assign w8238 = w1245 & ~w1377;
assign w8239 = ~w1371 & ~w1253;
assign w8240 = ~w1271 & w1266;
assign w8241 = ~pi01 & pi51;
assign w8242 = ~w1397 & ~w1396;
assign w8243 = ~pi00 & pi51;
assign w8244 = ~w1262 & w1404;
assign w8245 = w1303 & ~w1279;
assign w8246 = ~w1309 & w1412;
assign w8247 = w1309 & ~w1412;
assign w8248 = ~pi05 & pi47;
assign w8249 = ~w1431 & ~w1430;
assign w8250 = ~pi03 & pi49;
assign w8251 = ~w1437 & ~w1436;
assign w8252 = ~pi11 & pi41;
assign w8253 = ~w1462 & ~w1461;
assign w8254 = ~pi09 & pi43;
assign w8255 = ~w1468 & ~w1467;
assign w8256 = ~pi17 & pi35;
assign w8257 = ~w1483 & ~w1482;
assign w8258 = ~pi15 & pi37;
assign w8259 = ~w1489 & ~w1488;
assign w8260 = ~w1513 & ~w1387;
assign w8261 = ~w1408 & ~w1407;
assign w8262 = ~pi00 & ~pi53;
assign w8263 = ~w1394 & ~w1550;
assign w8264 = ~w1446 & ~w1422;
assign w8265 = ~pi06 & pi47;
assign w8266 = ~w1579 & ~w1578;
assign w8267 = ~pi04 & pi49;
assign w8268 = ~w1588 & ~w1587;
assign w8269 = ~pi18 & pi35;
assign w8270 = ~w1606 & ~w1605;
assign w8271 = ~pi16 & pi37;
assign w8272 = ~w1612 & ~w1611;
assign w8273 = ~pi10 & pi43;
assign w8274 = ~w1643 & ~w1642;
assign w8275 = ~pi12 & pi41;
assign w8276 = ~w1652 & ~w1651;
assign w8277 = w1522 & w1679;
assign w8278 = ~w1522 & ~w1679;
assign w8279 = ~pi00 & pi55;
assign w8280 = pi00 & ~pi55;
assign w8281 = ~pi01 & pi53;
assign w8282 = ~w1701 & ~w1700;
assign w8283 = w1709 & pi51;
assign w8284 = ~w1709 & ~pi51;
assign w8285 = ~w1582 & ~w1591;
assign w8286 = ~w1646 & ~w1655;
assign w8287 = ~pi07 & pi47;
assign w8288 = ~w1749 & ~w1748;
assign w8289 = ~pi05 & pi49;
assign w8290 = ~w1758 & ~w1757;
assign w8291 = ~pi17 & pi37;
assign w8292 = ~w1776 & ~w1775;
assign w8293 = ~pi19 & pi35;
assign w8294 = ~w1782 & ~w1781;
assign w8295 = ~pi11 & pi43;
assign w8296 = ~w1810 & ~w1809;
assign w8297 = ~pi13 & pi41;
assign w8298 = ~w1819 & ~w1818;
assign w8299 = w1679 & w1847;
assign w8300 = w1692 & ~w1722;
assign w8301 = ~pi02 & pi53;
assign w8302 = ~w1874 & ~w1873;
assign w8303 = ~w1813 & ~w1822;
assign w8304 = ~w1752 & ~w1761;
assign w8305 = ~pi06 & pi49;
assign w8306 = ~w1916 & ~w1915;
assign w8307 = ~pi08 & pi47;
assign w8308 = ~w1925 & ~w1924;
assign w8309 = ~pi20 & pi35;
assign w8310 = ~w1943 & ~w1942;
assign w8311 = ~pi18 & pi37;
assign w8312 = ~w1949 & ~w1948;
assign w8313 = ~pi12 & pi43;
assign w8314 = ~w1977 & ~w1976;
assign w8315 = ~pi14 & pi41;
assign w8316 = ~w1986 & ~w1985;
assign w8317 = ~w2372 & w2014;
assign w8318 = ~w2011 & ~w2010;
assign w8319 = ~w1855 & ~w1854;
assign w8320 = w1891 & ~w1888;
assign w8321 = ~w1897 & w2023;
assign w8322 = w1897 & ~w2023;
assign w8323 = ~pi00 & ~pi57;
assign w8324 = pi00 & pi57;
assign w8325 = w1877 & w2035;
assign w8326 = ~w1877 & ~w2035;
assign w8327 = ~pi01 & pi55;
assign w8328 = ~w2059 & ~w2058;
assign w8329 = ~w1980 & ~w1989;
assign w8330 = ~w1919 & ~w1928;
assign w8331 = ~pi07 & pi49;
assign w8332 = ~w2108 & ~w2107;
assign w8333 = ~pi13 & pi43;
assign w8334 = ~w2141 & ~w2140;
assign w8335 = w2155 & pi35;
assign w8336 = ~w2155 & ~pi35;
assign w8337 = ~pi19 & pi37;
assign w8338 = ~w2161 & ~w2160;
assign w8339 = w2193 & ~w2010;
assign w8340 = w2193 & w8318;
assign w8341 = w2075 & ~w2072;
assign w8342 = ~pi02 & pi55;
assign w8343 = ~w2231 & ~w2230;
assign w8344 = w2123 & ~w2124;
assign w8345 = ~w2158 & ~w2171;
assign w8346 = ~pi14 & pi43;
assign w8347 = ~w2314 & ~w2313;
assign w8348 = ~w2027 & w2021;
assign w8349 = w2248 & ~w2245;
assign w8350 = w2253 & ~w2395;
assign w8351 = ~w2253 & w2395;
assign w8352 = w2408 & pi57;
assign w8353 = ~w2408 & ~pi57;
assign w8354 = w2235 & ~w2411;
assign w8355 = ~pi55 & pi03;
assign w8356 = ~w2427 & ~w2429;
assign w8357 = ~pi05 & pi53;
assign w8358 = pi06 & pi53;
assign w8359 = w2438 & ~w2440;
assign w8360 = ~pi47 & pi11;
assign w8361 = ~w2471 & ~w2472;
assign w8362 = ~pi09 & pi49;
assign w8363 = ~pi49 & pi09;
assign w8364 = ~w2480 & ~w2482;
assign w8365 = ~pi41 & pi17;
assign w8366 = ~w2507 & ~w2508;
assign w8367 = ~pi15 & pi43;
assign w8368 = pi16 & pi43;
assign w8369 = w2517 & ~w2519;
assign w8370 = ~pi37 & pi21;
assign w8371 = ~w2528 & ~w2529;
assign w8372 = ~pi35 & pi23;
assign w8373 = ~w2534 & ~w2535;
assign w8374 = w2569 & w2572;
assign w8375 = w2569 & ~w8018;
assign w8376 = w2447 & ~w2404;
assign w8377 = pi00 & pi59;
assign w8378 = w2390 & w9091;
assign w8379 = ~w2590 & ~w2585;
assign w8380 = ~w2453 & w2596;
assign w8381 = w2453 & ~w2596;
assign w8382 = w2413 & ~w2414;
assign w8383 = w2609 & pi57;
assign w8384 = ~w2609 & ~pi57;
assign w8385 = ~w2432 & ~w2441;
assign w8386 = ~pi55 & pi04;
assign w8387 = ~w2626 & ~w2627;
assign w8388 = ~pi06 & pi53;
assign w8389 = pi07 & pi53;
assign w8390 = w2636 & ~w2638;
assign w8391 = ~w2498 & w2550;
assign w8392 = ~w2511 & ~w2520;
assign w8393 = ~w2475 & ~w2485;
assign w8394 = ~pi49 & pi10;
assign w8395 = ~w2671 & ~w2672;
assign w8396 = ~pi12 & pi47;
assign w8397 = pi13 & pi47;
assign w8398 = w2681 & ~w2683;
assign w8399 = ~pi22 & pi37;
assign w8400 = ~w2697 & ~w2696;
assign w8401 = ~pi24 & pi35;
assign w8402 = ~w2703 & ~w2702;
assign w8403 = pi41 & pi16;
assign w8404 = ~w2730 & ~w2731;
assign w8405 = ~pi18 & pi41;
assign w8406 = pi19 & pi41;
assign w8407 = w2740 & ~w2742;
assign w8408 = ~w2758 & ~w2768;
assign w8409 = w2453 & w2595;
assign w8410 = ~w2771 & ~w2770;
assign w8411 = w2615 & ~w2616;
assign w8412 = w2661 & ~w2660;
assign w8413 = w2783 & pi57;
assign w8414 = ~w2783 & ~pi57;
assign w8415 = ~w2630 & ~w2639;
assign w8416 = ~pi55 & pi05;
assign w8417 = ~w2800 & ~w2801;
assign w8418 = ~pi07 & pi53;
assign w8419 = pi08 & pi53;
assign w8420 = w2810 & ~w2812;
assign w8421 = ~w2675 & ~w2684;
assign w8422 = ~w2734 & ~w2743;
assign w8423 = ~pi49 & pi11;
assign w8424 = ~w2843 & ~w2844;
assign w8425 = ~pi13 & pi47;
assign w8426 = pi14 & pi47;
assign w8427 = w2853 & ~w2855;
assign w8428 = ~pi25 & pi35;
assign w8429 = ~w2871 & ~w2870;
assign w8430 = ~pi23 & pi37;
assign w8431 = ~w2877 & ~w2876;
assign w8432 = ~pi19 & pi41;
assign w8433 = ~w2905 & ~w2904;
assign w8434 = ~pi17 & pi43;
assign w8435 = ~w2914 & ~w2913;
assign w8436 = w2935 & pi59;
assign w8437 = ~w2935 & ~pi59;
assign w8438 = ~pi00 & pi59;
assign w8439 = ~w2590 & w2942;
assign w8440 = ~w2645 & ~w2605;
assign w8441 = ~w2652 & w2950;
assign w8442 = w2652 & ~w2950;
assign w8443 = w2568 & w2761;
assign w8444 = w2968 & w2964;
assign w8445 = ~w2968 & ~w2964;
assign w8446 = ~w2946 & ~w2945;
assign w8447 = w2983 & pi61;
assign w8448 = ~w2983 & ~pi61;
assign w8449 = w2988 & pi59;
assign w8450 = ~w2988 & ~pi59;
assign w8451 = ~pi00 & pi61;
assign w8452 = ~w2933 & ~w2995;
assign w8453 = ~w2819 & ~w2780;
assign w8454 = w2789 & ~w2790;
assign w8455 = w2833 & ~w2832;
assign w8456 = w3014 & pi57;
assign w8457 = ~w3014 & ~pi57;
assign w8458 = ~w2804 & ~w2813;
assign w8459 = ~pi08 & pi53;
assign w8460 = ~w3032 & ~w3031;
assign w8461 = ~pi06 & pi55;
assign w8462 = ~w3041 & ~w3040;
assign w8463 = ~w2908 & ~w2917;
assign w8464 = ~w2847 & ~w2856;
assign w8465 = ~pi12 & pi49;
assign w8466 = ~w3075 & ~w3074;
assign w8467 = ~pi14 & pi47;
assign w8468 = ~w3084 & ~w3083;
assign w8469 = ~pi24 & pi37;
assign w8470 = ~w3102 & ~w3101;
assign w8471 = ~pi26 & pi35;
assign w8472 = ~w3108 & ~w3107;
assign w8473 = ~pi20 & pi41;
assign w8474 = ~w3136 & ~w3135;
assign w8475 = ~pi18 & pi43;
assign w8476 = ~w3145 & ~w3144;
assign w8477 = w2569 & w2369;
assign w8478 = ~w3169 & ~w2383;
assign w8479 = ~pi00 & pi63;
assign w8480 = pi00 & ~pi63;
assign w8481 = w3191 & pi61;
assign w8482 = ~w3191 & ~pi61;
assign w8483 = w3199 & pi59;
assign w8484 = ~w3199 & ~pi59;
assign w8485 = w3050 & ~w3011;
assign w8486 = w3056 & ~w3218;
assign w8487 = ~w3056 & w3218;
assign w8488 = w3020 & ~w3021;
assign w8489 = w3064 & ~w3063;
assign w8490 = w3230 & pi57;
assign w8491 = ~w3230 & ~pi57;
assign w8492 = ~w3035 & ~w3044;
assign w8493 = ~pi09 & pi53;
assign w8494 = ~w3248 & ~w3247;
assign w8495 = ~pi07 & pi55;
assign w8496 = ~w3257 & ~w3256;
assign w8497 = ~w3078 & ~w3087;
assign w8498 = ~w3139 & ~w3148;
assign w8499 = ~pi13 & pi49;
assign w8500 = ~w3291 & ~w3290;
assign w8501 = ~pi15 & pi47;
assign w8502 = ~w3300 & ~w3299;
assign w8503 = ~pi25 & pi37;
assign w8504 = ~w3318 & ~w3317;
assign w8505 = ~pi27 & pi35;
assign w8506 = ~w3324 & ~w3323;
assign w8507 = ~pi21 & pi41;
assign w8508 = ~w3352 & ~w3351;
assign w8509 = ~pi19 & pi43;
assign w8510 = ~w3361 & ~w3360;
assign w8511 = ~w3167 & ~w3386;
assign w8512 = w3167 & w3386;
assign w8513 = w3379 & ~w3180;
assign w8514 = w3202 & ~w3195;
assign w8515 = w3398 & pi59;
assign w8516 = ~w3398 & ~pi59;
assign w8517 = w3406 & pi63;
assign w8518 = ~w3406 & ~pi63;
assign w8519 = w3411 & pi61;
assign w8520 = ~w3411 & ~pi61;
assign w8521 = ~w3208 & ~w3206;
assign w8522 = w3266 & ~w3227;
assign w8523 = w3272 & ~w3431;
assign w8524 = ~w3272 & w3431;
assign w8525 = w3280 & ~w3279;
assign w8526 = w3237 & ~w3236;
assign w8527 = w3443 & pi57;
assign w8528 = ~w3443 & ~pi57;
assign w8529 = ~w3251 & ~w3260;
assign w8530 = ~pi10 & pi53;
assign w8531 = ~w3461 & ~w3460;
assign w8532 = ~pi08 & pi55;
assign w8533 = ~w3470 & ~w3469;
assign w8534 = ~w3294 & ~w3303;
assign w8535 = ~w3355 & ~w3364;
assign w8536 = ~pi16 & pi47;
assign w8537 = ~w3504 & ~w3503;
assign w8538 = ~pi14 & pi49;
assign w8539 = ~w3513 & ~w3512;
assign w8540 = ~pi28 & pi35;
assign w8541 = ~w3537 & ~w3536;
assign w8542 = ~pi26 & pi37;
assign w8543 = ~w3543 & ~w3542;
assign w8544 = ~pi22 & pi41;
assign w8545 = ~w3565 & ~w3564;
assign w8546 = ~pi20 & pi43;
assign w8547 = ~w3574 & ~w3573;
assign w8548 = ~w3607 & w3598;
assign w8549 = w3607 & ~w3598;
assign w8550 = ~w3384 & ~w3597;
assign w8551 = ~w2382 & ~w3611;
assign w8552 = ~w3616 & ~w3611;
assign w8553 = ~w3592 & ~w3393;
assign w8554 = ~w3401 & ~w3415;
assign w8555 = w3628 & pi59;
assign w8556 = ~w3628 & ~pi59;
assign w8557 = w3633 & pi63;
assign w8558 = ~w3633 & ~pi63;
assign w8559 = w3638 & pi61;
assign w8560 = ~w3638 & ~pi61;
assign w8561 = w3479 & ~w3439;
assign w8562 = w3485 & w3657;
assign w8563 = ~w3485 & ~w3657;
assign w8564 = w3493 & ~w3492;
assign w8565 = w3449 & ~w3450;
assign w8566 = w3669 & pi57;
assign w8567 = ~w3669 & ~pi57;
assign w8568 = ~w3464 & ~w3473;
assign w8569 = ~pi11 & pi53;
assign w8570 = ~w3687 & ~w3686;
assign w8571 = ~pi09 & pi55;
assign w8572 = ~w3696 & ~w3695;
assign w8573 = ~w3507 & ~w3516;
assign w8574 = ~w3568 & ~w3577;
assign w8575 = ~pi17 & pi47;
assign w8576 = ~w3730 & ~w3729;
assign w8577 = ~pi15 & pi49;
assign w8578 = ~w3739 & ~w3738;
assign w8579 = ~pi21 & pi43;
assign w8580 = ~w3792 & ~w3791;
assign w8581 = ~pi23 & pi41;
assign w8582 = ~w3801 & ~w3800;
assign w8583 = ~w3596 & w3825;
assign w8584 = w3596 & ~w3825;
assign w8585 = w3819 & ~w3623;
assign w8586 = ~w3631 & ~w3642;
assign w8587 = w3837 & pi59;
assign w8588 = ~w3837 & ~pi59;
assign w8589 = ~w3705 & ~w3666;
assign w8590 = ~w3711 & w3866;
assign w8591 = w3711 & ~w3866;
assign w8592 = w3751 & ~w3752;
assign w8593 = w3719 & ~w3718;
assign w8594 = w3676 & ~w3675;
assign w8595 = w3879 & pi57;
assign w8596 = ~w3879 & ~pi57;
assign w8597 = ~w3690 & ~w3699;
assign w8598 = ~pi12 & pi53;
assign w8599 = ~w3896 & ~w3895;
assign w8600 = ~pi10 & pi55;
assign w8601 = ~w3905 & ~w3904;
assign w8602 = ~w3733 & ~w3742;
assign w8603 = ~w3795 & ~w3804;
assign w8604 = ~pi18 & pi47;
assign w8605 = ~w3937 & ~w3936;
assign w8606 = ~pi16 & pi49;
assign w8607 = ~w3946 & ~w3945;
assign w8608 = ~w4021 & ~w3823;
assign w8609 = ~w4021 & w8020;
assign w8610 = ~w4015 & ~w3832;
assign w8611 = ~w3840 & ~w3851;
assign w8612 = w4035 & pi59;
assign w8613 = ~w4035 & ~pi59;
assign w8614 = w4071 & pi57;
assign w8615 = ~w4071 & ~pi57;
assign w8616 = ~w3899 & ~w3908;
assign w8617 = ~pi11 & pi55;
assign w8618 = ~w4088 & ~w4087;
assign w8619 = ~pi13 & pi53;
assign w8620 = ~w4097 & ~w4096;
assign w8621 = w3926 & ~w3925;
assign w8622 = ~w3940 & ~w3949;
assign w8623 = ~pi19 & pi47;
assign w8624 = ~w4136 & ~w4135;
assign w8625 = ~pi17 & pi49;
assign w8626 = ~w4145 & ~w4144;
assign w8627 = ~pi23 & pi43;
assign w8628 = ~w4191 & ~w4190;
assign w8629 = ~pi25 & pi41;
assign w8630 = ~w4200 & ~w4199;
assign w8631 = w4227 & ~w1680;
assign w8632 = w4228 & ~w4239;
assign w8633 = w7892 & w4224;
assign w8634 = (w4224 & w7892) | (w4224 & ~w4228) | (w7892 & ~w4228);
assign w8635 = w4068 & w4245;
assign w8636 = ~w4058 & w4065;
assign w8637 = ~w4058 & w7650;
assign w8638 = ~w4038 & ~w4049;
assign w8639 = w4255 & pi59;
assign w8640 = ~w4255 & ~pi59;
assign w8641 = ~w4091 & ~w4100;
assign w8642 = w4300 & pi51;
assign w8643 = ~w4300 & ~pi51;
assign w8644 = ~pi14 & pi53;
assign w8645 = ~w4306 & ~w4305;
assign w8646 = ~pi12 & pi55;
assign w8647 = ~w4312 & ~w4311;
assign w8648 = w4151 & ~w4124;
assign w8649 = ~w4139 & ~w4148;
assign w8650 = ~w4194 & ~w4203;
assign w8651 = w4029 & ~w4030;
assign w8652 = w4222 & ~w4223;
assign w8653 = ~w4434 & ~w8633;
assign w8654 = (w8022 & w8021) | (w8022 & w4228) | (w8021 & w4228);
assign w8655 = ~w4249 & w4244;
assign w8656 = ~w4425 & ~w4439;
assign w8657 = ~w4258 & ~w4269;
assign w8658 = w4443 & pi59;
assign w8659 = ~w4443 & ~pi59;
assign w8660 = w4448 & pi63;
assign w8661 = ~w4448 & ~pi63;
assign w8662 = w4453 & pi61;
assign w8663 = ~w4453 & ~pi61;
assign w8664 = w4329 & ~w4326;
assign w8665 = ~w4321 & ~w4297;
assign w8666 = w4303 & ~w4316;
assign w8667 = w4480 & pi57;
assign w8668 = ~w4480 & ~pi57;
assign w8669 = ~pi15 & pi53;
assign w8670 = ~w4493 & ~w4492;
assign w8671 = ~pi13 & pi55;
assign w8672 = ~w4502 & ~w4501;
assign w8673 = ~pi19 & pi49;
assign w8674 = ~w4534 & ~w4533;
assign w8675 = ~pi21 & pi47;
assign w8676 = ~w4543 & ~w4542;
assign w8677 = ~pi27 & pi41;
assign w8678 = ~w4560 & ~w4559;
assign w8679 = ~pi25 & pi43;
assign w8680 = ~w4566 & ~w4565;
assign w8681 = ~pi31 & ~pi37;
assign w8682 = pi37 & pi31;
assign w8683 = ~pi29 & pi39;
assign w8684 = ~w4581 & ~w4580;
assign w8685 = ~w4626 & ~w4431;
assign w8686 = ~w4626 & w8023;
assign w8687 = ~w4468 & ~w4466;
assign w8688 = w4483 & w4478;
assign w8689 = w4648 & pi57;
assign w8690 = ~w4648 & ~pi57;
assign w8691 = ~w4496 & ~w4505;
assign w8692 = ~pi14 & pi55;
assign w8693 = ~w4663 & ~w4662;
assign w8694 = ~pi16 & pi53;
assign w8695 = ~w4669 & ~w4668;
assign w8696 = w4549 & ~w4522;
assign w8697 = ~pi26 & pi43;
assign w8698 = ~w4703 & ~w4702;
assign w8699 = ~pi28 & pi41;
assign w8700 = ~w4712 & ~w4711;
assign w8701 = ~w4537 & ~w4546;
assign w8702 = ~pi20 & pi49;
assign w8703 = ~w4738 & ~w4737;
assign w8704 = ~pi22 & pi47;
assign w8705 = ~w4747 & ~w4746;
assign w8706 = ~w4446 & ~w4457;
assign w8707 = w4769 & pi59;
assign w8708 = ~w4769 & ~pi59;
assign w8709 = w4774 & pi63;
assign w8710 = ~w4774 & ~pi63;
assign w8711 = w4779 & pi61;
assign w8712 = ~w4779 & ~pi61;
assign w8713 = ~w4475 & w4794;
assign w8714 = w4475 & ~w4794;
assign w8715 = ~w4820 & w4810;
assign w8716 = w4820 & ~w4810;
assign w8717 = ~w4688 & ~w4762;
assign w8718 = w4727 & ~w4726;
assign w8719 = w4839 & pi57;
assign w8720 = ~w4839 & ~pi57;
assign w8721 = w4673 & ~w4842;
assign w8722 = ~pi17 & pi53;
assign w8723 = ~w4856 & ~w4855;
assign w8724 = ~pi15 & pi55;
assign w8725 = ~w4865 & ~w4864;
assign w8726 = ~pi29 & pi41;
assign w8727 = ~w4880 & ~w4879;
assign w8728 = ~pi27 & pi43;
assign w8729 = ~w4886 & ~w4885;
assign w8730 = ~pi31 & pi39;
assign w8731 = ~w4741 & ~w4750;
assign w8732 = ~w4706 & ~w4715;
assign w8733 = ~pi23 & pi47;
assign w8734 = ~w4919 & ~w4918;
assign w8735 = ~pi21 & pi49;
assign w8736 = ~w4928 & ~w4927;
assign w8737 = w4685 & ~w4683;
assign w8738 = ~w4772 & ~w4783;
assign w8739 = w4954 & pi59;
assign w8740 = ~w4954 & ~pi59;
assign w8741 = w4959 & pi63;
assign w8742 = ~w4959 & ~pi63;
assign w8743 = w4964 & pi61;
assign w8744 = ~w4964 & ~pi61;
assign w8745 = ~w4239 & w4991;
assign w8746 = ~w4998 & w5002;
assign w8747 = ~w4979 & ~w4977;
assign w8748 = ~w4957 & ~w4968;
assign w8749 = w5017 & pi59;
assign w8750 = ~w5017 & ~pi59;
assign w8751 = w5053 & pi41;
assign w8752 = ~w5053 & ~pi41;
assign w8753 = w5060 & pi43;
assign w8754 = ~w5060 & ~pi43;
assign w8755 = ~w4922 & ~w4931;
assign w8756 = ~pi24 & pi47;
assign w8757 = ~w5083 & ~w5082;
assign w8758 = ~pi22 & pi49;
assign w8759 = ~w5092 & ~w5091;
assign w8760 = w4844 & ~w4845;
assign w8761 = w4907 & ~w4908;
assign w8762 = w5115 & pi57;
assign w8763 = ~w5115 & ~pi57;
assign w8764 = ~w4859 & ~w4868;
assign w8765 = ~pi18 & pi53;
assign w8766 = ~w5132 & ~w5131;
assign w8767 = ~pi16 & pi55;
assign w8768 = ~w5141 & ~w5140;
assign w8769 = ~w5165 & w4996;
assign w8770 = ~w5165 & w8024;
assign w8771 = ~w5020 & ~w5031;
assign w8772 = w5177 & pi59;
assign w8773 = ~w5177 & ~pi59;
assign w8774 = w5072 & ~w5071;
assign w8775 = w5217 & pi57;
assign w8776 = ~w5217 & ~pi57;
assign w8777 = ~w5135 & ~w5144;
assign w8778 = ~pi19 & pi53;
assign w8779 = ~w5235 & ~w5234;
assign w8780 = ~pi17 & pi55;
assign w8781 = ~w5244 & ~w5243;
assign w8782 = ~w5086 & ~w5095;
assign w8783 = w5263 & pi43;
assign w8784 = ~w5263 & ~pi43;
assign w8785 = ~pi31 & pi41;
assign w8786 = ~pi23 & pi49;
assign w8787 = ~w5283 & ~w5282;
assign w8788 = ~pi25 & pi47;
assign w8789 = ~w5292 & ~w5291;
assign w8790 = w5164 & ~w5163;
assign w8791 = ~w5320 & ~w5331;
assign w8792 = w5256 & ~w5305;
assign w8793 = w5259 & ~w5260;
assign w8794 = w5223 & ~w5224;
assign w8795 = w5346 & pi57;
assign w8796 = ~w5346 & ~pi57;
assign w8797 = ~w5238 & ~w5247;
assign w8798 = ~pi20 & pi53;
assign w8799 = ~w5364 & ~w5363;
assign w8800 = ~pi18 & pi55;
assign w8801 = ~w5373 & ~w5372;
assign w8802 = ~w5286 & ~w5295;
assign w8803 = w5395 & pi45;
assign w8804 = ~w5395 & ~pi45;
assign w8805 = ~pi24 & pi49;
assign w8806 = ~w5401 & ~w5400;
assign w8807 = ~pi26 & pi47;
assign w8808 = ~w5407 & ~w5406;
assign w8809 = ~pi30 & ~w355;
assign w8810 = ~w5180 & ~w5191;
assign w8811 = w5449 & pi59;
assign w8812 = ~w5449 & ~pi59;
assign w8813 = w5454 & pi63;
assign w8814 = ~w5454 & ~pi63;
assign w8815 = w5459 & pi61;
assign w8816 = ~w5459 & ~pi61;
assign w8817 = w5253 & ~w5214;
assign w8818 = ~w5452 & ~w5463;
assign w8819 = w5518 & pi59;
assign w8820 = ~w5518 & ~pi59;
assign w8821 = w5523 & pi63;
assign w8822 = ~w5523 & ~pi63;
assign w8823 = w5528 & pi61;
assign w8824 = ~w5528 & ~pi61;
assign w8825 = w5352 & ~w5353;
assign w8826 = w5558 & pi57;
assign w8827 = ~w5558 & ~pi57;
assign w8828 = ~w5367 & ~w5376;
assign w8829 = w5603 & pi45;
assign w8830 = ~w5603 & ~pi45;
assign w8831 = w5165 & w4809;
assign w8832 = w7920 & ~w5496;
assign w8833 = (~w5496 & w7920) | (~w5496 & w5656) | (w7920 & w5656);
assign w8834 = ~w5521 & ~w5532;
assign w8835 = w5673 & pi59;
assign w8836 = ~w5673 & ~pi59;
assign w8837 = w5597 & ~w5634;
assign w8838 = ~w5606 & ~w5621;
assign w8839 = w5709 & pi45;
assign w8840 = ~w5709 & ~pi45;
assign w8841 = w5564 & ~w5565;
assign w8842 = ~w5676 & ~w5687;
assign w8843 = w5819 & pi59;
assign w8844 = ~w5819 & ~pi59;
assign w8845 = ~pi31 & pi45;
assign w8846 = ~w5936 & ~w5801;
assign w8847 = ~w5822 & ~w5833;
assign w8848 = w5968 & pi59;
assign w8849 = ~w5968 & ~pi59;
assign w8850 = w6045 & pi49;
assign w8851 = ~w6045 & ~pi49;
assign w8852 = w6051 & pi47;
assign w8853 = ~w6051 & ~pi47;
assign w8854 = w5931 & ~w6086;
assign w8855 = ~w5938 & w8791;
assign w8856 = ~w5993 & ~w5991;
assign w8857 = ~pi31 & pi47;
assign w8858 = ~w5971 & ~w5982;
assign w8859 = w6175 & pi59;
assign w8860 = ~w6175 & ~pi59;
assign w8861 = w6214 & w5930;
assign w8862 = ~w6178 & ~w6189;
assign w8863 = w6234 & pi59;
assign w8864 = ~w6234 & ~pi59;
assign w8865 = w6266 & pi57;
assign w8866 = ~w6266 & ~pi57;
assign w8867 = w6306 & pi49;
assign w8868 = ~w6306 & ~pi49;
assign w8869 = ~w6056 & ~w6309;
assign w8870 = w6097 & ~w6098;
assign w8871 = ~w6259 & ~w6257;
assign w8872 = w6321 & w6344;
assign w8873 = ~w6321 & ~w6344;
assign w8874 = ~w6237 & ~w6248;
assign w8875 = w6353 & pi59;
assign w8876 = ~w6353 & ~pi59;
assign w8877 = w6302 & w6162;
assign w8878 = ~pi31 & pi49;
assign w8879 = ~w6309 & w6437;
assign w8880 = w5648 & w5653;
assign w8881 = ~w6356 & ~w6367;
assign w8882 = w6488 & pi59;
assign w8883 = ~w6488 & ~pi59;
assign w8884 = ~w5932 & w5936;
assign w8885 = ~pi31 & pi51;
assign w8886 = w6620 & pi57;
assign w8887 = ~w6620 & ~pi57;
assign w8888 = ~w6491 & ~w6502;
assign w8889 = w6636 & pi59;
assign w8890 = ~w6636 & ~pi59;
assign w8891 = w6696 & pi55;
assign w8892 = ~w6696 & ~pi55;
assign w8893 = w6702 & pi53;
assign w8894 = ~w6702 & ~pi53;
assign w8895 = w6711 & pi57;
assign w8896 = ~w6711 & ~pi57;
assign w8897 = w6617 & ~w6624;
assign w8898 = w6727 & pi59;
assign w8899 = ~w6727 & ~pi59;
assign w8900 = ~w6757 & ~w6659;
assign w8901 = w6677 & ~w6767;
assign w8902 = ~w6677 & ~w6771;
assign w8903 = w6677 & ~w6775;
assign w8904 = w5945 & ~w4990;
assign w8905 = (~w6782 & w5333) | (~w6782 & w8996) | (w5333 & w8996);
assign w8906 = ~w6786 & w5328;
assign w8907 = w6798 & pi55;
assign w8908 = ~w6798 & ~pi55;
assign w8909 = ~pi31 & pi53;
assign w8910 = w6810 & pi57;
assign w8911 = ~w6810 & ~pi57;
assign w8912 = w6708 & ~w6716;
assign w8913 = ~w6730 & ~w6739;
assign w8914 = w6826 & pi59;
assign w8915 = ~w6826 & ~pi59;
assign w8916 = w6724 & w6748;
assign w8917 = ~w6724 & ~w6748;
assign w8918 = w6694 & ~w6759;
assign w8919 = w6765 & w6868;
assign w8920 = ~w6765 & ~w6868;
assign w8921 = w6685 & w6873;
assign w8922 = ~w6685 & ~w6877;
assign w8923 = ~w6857 & ~w6858;
assign w8924 = ~w6808 & ~w6815;
assign w8925 = w6900 & pi55;
assign w8926 = ~w6900 & ~pi55;
assign w8927 = w6905 & pi57;
assign w8928 = ~w6905 & ~pi57;
assign w8929 = ~w6829 & ~w6840;
assign w8930 = w6920 & pi59;
assign w8931 = ~w6920 & ~pi59;
assign w8932 = w6925 & pi63;
assign w8933 = ~w6925 & ~pi63;
assign w8934 = w6930 & pi61;
assign w8935 = ~w6930 & ~pi61;
assign w8936 = w6823 & w6849;
assign w8937 = ~w6823 & ~w6849;
assign w8938 = w6903 & ~w6909;
assign w8939 = w6972 & pi57;
assign w8940 = ~w6972 & ~pi57;
assign w8941 = ~pi31 & pi55;
assign w8942 = ~w6923 & ~w6934;
assign w8943 = w6991 & pi59;
assign w8944 = ~w6991 & ~pi59;
assign w8945 = w6996 & pi63;
assign w8946 = ~w6996 & ~pi63;
assign w8947 = w7001 & pi61;
assign w8948 = ~w7001 & ~pi61;
assign w8949 = w6917 & w6943;
assign w8950 = ~w4067 & w4244;
assign w8951 = ~w4247 & ~w4249;
assign w8952 = w4432 & w4223;
assign w8953 = w6895 & w7830;
assign w8954 = w7831 & ~w7330;
assign w8955 = (~w7330 & w7831) | (~w7330 & ~w6895) | (w7831 & ~w6895);
assign w8956 = w7384 & w7388;
assign w8957 = (w6962 & w6887) | (w6962 & w8997) | (w6887 & w8997);
assign w8958 = w6962 & ~w6894;
assign w8959 = w6967 & ~w6962;
assign w8960 = w6967 & ~w7962;
assign w8961 = ~w6917 & ~w6943;
assign w8962 = ~w6866 & ~w6959;
assign w8963 = ~w7064 & ~w7074;
assign w8964 = w7057 & w7083;
assign w8965 = ~w7057 & ~w7083;
assign w8966 = w6464 & w7166;
assign w8967 = ~w7828 & w7184;
assign w8968 = w7118 & w7144;
assign w8969 = ~w7118 & ~w7144;
assign w8970 = ~w7287 & w7289;
assign w8971 = w7040 & w7366;
assign w8972 = pi05 & pi45;
assign w8973 = ~pi05 & ~pi45;
assign w8974 = pi11 & pi39;
assign w8975 = ~pi11 & ~pi39;
assign w8976 = ~pi06 & ~pi45;
assign w8977 = pi12 & pi39;
assign w8978 = ~pi12 & ~pi39;
assign w8979 = pi08 & pi45;
assign w8980 = ~pi08 & ~pi45;
assign w8981 = pi14 & pi39;
assign w8982 = ~pi14 & ~pi39;
assign w8983 = ~w2080 & ~w2197;
assign w8984 = w2080 & w2197;
assign w8985 = pi23 & pi35;
assign w8986 = ~pi23 & ~pi35;
assign w8987 = ~pi21 & ~pi37;
assign w8988 = w5319 & w5164;
assign w8989 = w4797 & ~w4827;
assign w8990 = ~w4797 & w4827;
assign w8991 = ~w3617 & w6782;
assign w8992 = w7828 & ~w7285;
assign w8993 = ~w7283 & ~w8009;
assign w8994 = ~w7283 & ~w8010;
assign w8995 = w6464 & w4815;
assign w8996 = ~w6785 & ~w6782;
assign w8997 = w6792 & w6962;
assign w8998 = pi03 & pi47;
assign w8999 = pi01 & pi49;
assign w9000 = pi09 & pi41;
assign w9001 = pi07 & pi43;
assign w9002 = pi04 & pi47;
assign w9003 = pi02 & pi49;
assign w9004 = pi10 & pi41;
assign w9005 = pi08 & pi43;
assign w9006 = pi06 & pi47;
assign w9007 = pi04 & pi49;
assign w9008 = pi12 & pi41;
assign w9009 = pi10 & pi43;
assign w9010 = pi04 & pi55;
assign w9011 = ~pi53 & pi05;
assign w9012 = pi12 & pi47;
assign w9013 = pi10 & pi49;
assign w9014 = pi18 & pi41;
assign w9015 = pi41 & pi15;
assign w9016 = pi22 & pi37;
assign w9017 = pi24 & pi35;
assign w9018 = pi05 & pi55;
assign w9019 = ~pi53 & pi06;
assign w9020 = pi11 & pi49;
assign w9021 = ~pi47 & pi12;
assign w9022 = pi23 & pi37;
assign w9023 = pi25 & pi35;
assign w9024 = pi17 & pi43;
assign w9025 = ~pi41 & pi18;
assign w9026 = pi06 & pi55;
assign w9027 = ~pi53 & pi07;
assign w9028 = pi12 & pi49;
assign w9029 = ~pi47 & pi13;
assign w9030 = pi26 & pi35;
assign w9031 = pi24 & pi37;
assign w9032 = pi20 & pi41;
assign w9033 = pi18 & pi43;
assign w9034 = pi09 & pi53;
assign w9035 = pi07 & pi55;
assign w9036 = pi13 & pi49;
assign w9037 = pi15 & pi47;
assign w9038 = pi25 & pi37;
assign w9039 = pi27 & pi35;
assign w9040 = pi21 & pi41;
assign w9041 = pi19 & pi43;
assign w9042 = pi10 & pi53;
assign w9043 = pi08 & pi55;
assign w9044 = pi14 & pi49;
assign w9045 = pi16 & pi47;
assign w9046 = pi26 & pi37;
assign w9047 = pi28 & pi35;
assign w9048 = pi22 & pi41;
assign w9049 = pi20 & pi43;
assign w9050 = pi29 & pi35;
assign w9051 = pi27 & pi37;
assign w9052 = pi27 & pi43;
assign w9053 = pi29 & pi41;
assign w9054 = pi21 & pi49;
assign w9055 = pi23 & pi47;
assign w9056 = w4432 & w4224;
assign w9057 = pi30 & pi41;
assign w9058 = pi28 & pi43;
assign w9059 = pi24 & pi47;
assign w9060 = pi22 & pi49;
assign w9061 = w4991 & ~w4808;
assign w9062 = w4991 & w4815;
assign w9063 = pi25 & pi47;
assign w9064 = pi23 & pi49;
assign w9065 = pi19 & pi53;
assign w9066 = pi17 & pi55;
assign w9067 = pi20 & pi53;
assign w9068 = pi18 & pi55;
assign w9069 = pi24 & pi49;
assign w9070 = pi26 & pi47;
assign w9071 = ~w5332 & w5320;
assign w9072 = pi25 & pi49;
assign w9073 = pi27 & pi47;
assign w9074 = ~w6468 & ~w6466;
assign w9075 = ~w6468 & ~w3602;
assign w9076 = pi06 & pi45;
assign w9077 = pi21 & pi37;
assign w9078 = ~w684 & ~w687;
assign w9079 = (w2010 & ~w8318) | (w2010 & ~w2015) | (~w8318 & ~w2015);
assign w9080 = (~w2572 & w8018) | (~w2572 & ~w2383) | (w8018 & ~w2383);
assign w9081 = (w3173 & w2383) | (w3173 & ~w8019) | (w2383 & ~w8019);
assign w9082 = (~w3175 & ~w3169) | (~w3175 & w8478) | (~w3169 & w8478);
assign w9083 = (w3823 & ~w8020) | (w3823 & ~w3619) | (~w8020 & ~w3619);
assign w9084 = (w4431 & ~w8023) | (w4431 & ~w4630) | (~w8023 & ~w4630);
assign w9085 = (~w4996 & ~w8024) | (~w4996 & ~w8025) | (~w8024 & ~w8025);
assign w9086 = (w6081 & w6214) | (w6081 & w8861) | (w6214 & w8861);
assign w9087 = (~w5936 & ~w8884) | (~w5936 & ~w5656) | (~w8884 & ~w5656);
assign w9088 = (~w6093 & ~w8056) | (~w6093 & ~w5334) | (~w8056 & ~w5334);
assign w9089 = w8134 & pi01;
assign w9090 = w8220 & pi01;
assign w9091 = w8377 & pi01;
assign w9092 = (~w1520 & ~w7882) | (~w1520 & ~w1124) | (~w7882 & ~w1124);
assign w9093 = w5320 & ~w5333;
assign w9094 = (~w7043 & w7870) | (~w7043 & ~w6475) | (w7870 & ~w6475);
assign w9095 = (w8009 & w8010) | (w8009 & ~w6796) | (w8010 & ~w6796);
assign one = 1;
assign po00 = w0;
assign po01 = ~w5;
assign po02 = ~w21;
assign po03 = w47;
assign po04 = w80;
assign po05 = w116;
assign po06 = w157;
assign po07 = w211;
assign po08 = w272;
assign po09 = w344;
assign po10 = w424;
assign po11 = w517;
assign po12 = w602;
assign po13 = w689;
assign po14 = w779;
assign po15 = ~w888;
assign po16 = w1005;
assign po17 = w1128;
assign po18 = w1250;
assign po19 = ~w1384;
assign po20 = w1527;
assign po21 = ~w1683;
assign po22 = w1850;
assign po23 = w2018;
assign po24 = w2196;
assign po25 = w2386;
assign po26 = w2575;
assign po27 = ~w2767;
assign po28 = ~w2972;
assign po29 = w3178;
assign po30 = w3389;
assign po31 = w3610;
assign po32 = w3828;
assign po33 = w4025;
assign po34 = ~w4243;
assign po35 = w4438;
assign po36 = w4634;
assign po37 = w4824;
assign po38 = w5004;
assign po39 = w5168;
assign po40 = w5338;
assign po41 = w5503;
assign po42 = w5663;
assign po43 = w5808;
assign po44 = ~w5952;
assign po45 = w6090;
assign po46 = w6222;
assign po47 = ~w6343;
assign po48 = ~w6479;
assign po49 = ~w6584;
assign po50 = ~w6691;
assign po51 = ~w6781;
assign po52 = w6882;
assign po53 = w6969;
assign po54 = ~w7046;
assign po55 = w7110;
assign po56 = w7183;
assign po57 = ~w7243;
assign po58 = w7295;
assign po59 = w7333;
assign po60 = w7379;
assign po61 = ~w7414;
assign po62 = ~w7447;
assign po63 = ~w7454;
endmodule

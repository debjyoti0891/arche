module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371;
assign w0 = w244 & w136;
assign w1 = (w311 & w268) | (w311 & w199) | (w268 & w199);
assign w2 = (~pi004 & ~w281) | (~pi004 & w227) | (~w281 & w227);
assign w3 = ~pi022 & pi002;
assign w4 = w91 & w90;
assign w5 = (~pi041 & w264) | (~pi041 & w363) | (w264 & w363);
assign w6 = pi017 & pi073;
assign w7 = w249 & ~w245;
assign w8 = ~pi041 & pi042;
assign w9 = ~w111 & w350;
assign w10 = pi001 & pi099;
assign w11 = pi001 & w281;
assign w12 = pi073 & ~w47;
assign w13 = w139 & w17;
assign w14 = w53 & w100;
assign w15 = w311 & ~w268;
assign w16 = pi082 & pi089;
assign w17 = ~w299 & ~w239;
assign w18 = ~pi074 & pi081;
assign w19 = w261 & w7;
assign w20 = pi038 & pi043;
assign w21 = ~w336 & w349;
assign w22 = pi083 & ~pi087;
assign w23 = pi099 & ~w278;
assign w24 = ~w226 & ~w103;
assign w25 = (pi001 & w144) | (pi001 & w205) | (w144 & w205);
assign w26 = w77 & ~w85;
assign w27 = ~w59 & w35;
assign w28 = pi078 & ~w16;
assign w29 = w46 | ~w80;
assign w30 = ~w220 & w161;
assign w31 = pi084 & pi093;
assign w32 = ~pi019 & pi064;
assign w33 = ~w5 & w126;
assign w34 = pi079 & ~w31;
assign w35 = ~w351 & ~w72;
assign w36 = ~w111 & w70;
assign w37 = (~w355 & w29) | (~w355 & w258) | (w29 & w258);
assign w38 = pi056 & ~w94;
assign w39 = ~pi037 & ~pi110;
assign w40 = pi088 & ~pi032;
assign w41 = ~pi038 & ~pi043;
assign w42 = (~pi034 & ~w91) | (~pi034 & w182) | (~w91 & w182);
assign w43 = w63 & ~w279;
assign w44 = w166 & w67;
assign w45 = (~pi032 & ~w75) | (~pi032 & w40) | (~w75 & w40);
assign w46 = ~pi095 & ~w80;
assign w47 = ~w150 & ~w131;
assign w48 = ~pi066 & pi073;
assign w49 = w281 & w308;
assign w50 = w314 & w83;
assign w51 = ~w257 & w273;
assign w52 = ~pi037 & ~pi107;
assign w53 = ~w7 & ~w238;
assign w54 = ~w342 & ~w370;
assign w55 = pi033 & w63;
assign w56 = w325 & pi031;
assign w57 = pi095 & w337;
assign w58 = w311 & ~w41;
assign w59 = w144 & w355;
assign w60 = ~w111 & w266;
assign w61 = pi099 & ~w240;
assign w62 = w334 & ~w97;
assign w63 = pi073 & pi099;
assign w64 = ~w218 & w260;
assign w65 = ~pi058 & ~w73;
assign w66 = ~w165 & w251;
assign w67 = ~w323 & w45;
assign w68 = pi099 & ~w344;
assign w69 = ~w193 & ~w255;
assign w70 = ~w287 & ~w223;
assign w71 = ~w19 & w13;
assign w72 = pi002 & pi073;
assign w73 = ~pi070 & pi073;
assign w74 = ~w367 & w21;
assign w75 = pi041 & pi042;
assign w76 = ~w145 & ~w156;
assign w77 = pi000 & pi099;
assign w78 = w72 & w313;
assign w79 = pi099 & ~w250;
assign w80 = (pi002 & ~w288) | (pi002 & w3) | (~w288 & w3);
assign w81 = ~w111 & w338;
assign w82 = ~pi001 & w290;
assign w83 = pi027 & ~pi060;
assign w84 = ~w65 & w189;
assign w85 = pi034 & pi073;
assign w86 = ~w325 & ~pi031;
assign w87 = ~pi015 & pi037;
assign w88 = w334 & ~w152;
assign w89 = pi096 & w75;
assign w90 = pi056 & w94;
assign w91 = (pi073 & ~w280) | (pi073 & w85) | (~w280 & w85);
assign w92 = ~w39 & ~w225;
assign w93 = ~w180 & w339;
assign w94 = pi029 & pi034;
assign w95 = ~w12 & w116;
assign w96 = ~w111 & w107;
assign w97 = (~pi025 & ~w232) | (~pi025 & w222) | (~w232 & w222);
assign w98 = ~w264 & w179;
assign w99 = ~w286 & w77;
assign w100 = pi099 & pi104;
assign w101 = ~pi090 & w8;
assign w102 = ~w55 & ~w362;
assign w103 = pi007 & pi037;
assign w104 = ~w111 & w24;
assign w105 = ~w111 & w253;
assign w106 = ~w292 & ~w137;
assign w107 = ~w187 & ~w87;
assign w108 = ~w204 & ~w340;
assign w109 = pi032 & w75;
assign w110 = pi032 & w268;
assign w111 = w295 & w209;
assign w112 = pi053 & ~pi077;
assign w113 = pi094 & w8;
assign w114 = ~w25 & w0;
assign w115 = pi021 & w213;
assign w116 = pi002 & ~w167;
assign w117 = pi022 & ~pi073;
assign w118 = pi073 & w75;
assign w119 = ~pi044 & ~w117;
assign w120 = ~w186 & w364;
assign w121 = (~w290 & w2) | (~w290 & w318) | (w2 & w318);
assign w122 = pi059 & w293;
assign w123 = ~pi026 & ~pi024;
assign w124 = ~w18 & ~w135;
assign w125 = w312 & w78;
assign w126 = (w311 & w264) | (w311 & w195) | (w264 & w195);
assign w127 = w341 & w10;
assign w128 = pi099 & ~w177;
assign w129 = w32 & w53;
assign w130 = pi099 & ~w254;
assign w131 = ~pi074 & ~pi075;
assign w132 = w232 & w140;
assign w133 = pi020 & w91;
assign w134 = ~w309 & w283;
assign w135 = pi074 & ~pi081;
assign w136 = ~w49 & ~w82;
assign w137 = pi053 & w63;
assign w138 = pi058 & w73;
assign w139 = ~w111 & ~w50;
assign w140 = w188 & pi025;
assign w141 = pi099 & pi018;
assign w142 = ~pi010 & pi037;
assign w143 = (w77 & ~w91) | (w77 & w272) | (~w91 & w272);
assign w144 = pi005 & ~w2;
assign w145 = w315 & ~w303;
assign w146 = pi017 & ~pi027;
assign w147 = ~pi055 & w293;
assign w148 = (w77 & ~w91) | (w77 & w322) | (~w91 & w322);
assign w149 = ~w160 & ~w302;
assign w150 = pi074 & pi075;
assign w151 = pi019 & ~pi027;
assign w152 = pi026 & w232;
assign w153 = pi057 & w293;
assign w154 = w63 & ~w343;
assign w155 = pi020 & ~w91;
assign w156 = ~w43 & ~w122;
assign w157 = ~w264 & w211;
assign w158 = ~w234 & ~w157;
assign w159 = pi024 & pi025;
assign w160 = pi066 & w293;
assign w161 = w288 & w162;
assign w162 = pi002 & pi023;
assign w163 = ~w98 & ~w153;
assign w164 = pi072 & pi073;
assign w165 = (~pi001 & ~w328) | (~pi001 & w262) | (~w328 & w262);
assign w166 = ~w171 & ~w113;
assign w167 = pi056 & ~pi073;
assign w168 = ~pi002 & ~pi016;
assign w169 = pi000 & w91;
assign w170 = ~w158 & w58;
assign w171 = ~pi085 & w185;
assign w172 = w229 & w121;
assign w173 = pi073 & pi041;
assign w174 = ~pi057 & pi073;
assign w175 = ~w146 & ~w249;
assign w176 = ~w300 & w201;
assign w177 = ~w337 & ~w215;
assign w178 = pi033 & ~pi068;
assign w179 = w190 & w311;
assign w180 = (~pi054 & ~w73) | (~pi054 & w259) | (~w73 & w259);
assign w181 = ~w328 & ~w202;
assign w182 = ~pi056 & ~pi034;
assign w183 = pi043 & pi073;
assign w184 = w327 & w134;
assign w185 = pi041 & ~pi042;
assign w186 = ~pi072 & ~pi073;
assign w187 = ~pi037 & ~pi111;
assign w188 = pi026 & pi024;
assign w189 = w334 & ~w138;
assign w190 = pi073 & pi030;
assign w191 = ~w44 & w345;
assign w192 = ~w305 & w99;
assign w193 = pi067 & w63;
assign w194 = pi086 & pi032;
assign w195 = ~w173 & w311;
assign w196 = ~w271 & w88;
assign w197 = pi008 & w207;
assign w198 = ~pi041 & ~pi042;
assign w199 = pi032 & w311;
assign w200 = ~pi013 & pi037;
assign w201 = w77 & ~w228;
assign w202 = ~pi016 & ~pi073;
assign w203 = ~w124 & w57;
assign w204 = ~pi004 & ~w229;
assign w205 = w221 & w216;
assign w206 = ~w22 & ~w247;
assign w207 = pi003 & pi006;
assign w208 = ~w248 & w210;
assign w209 = ~pi027 & pi104;
assign w210 = pi099 & ~w48;
assign w211 = w190 & ~w20;
assign w212 = ~pi082 & ~pi084;
assign w213 = ~pi095 & ~pi018;
assign w214 = w159 & w235;
assign w215 = (w124 & w231) | (w124 & w115) | (w231 & w115);
assign w216 = pi095 & pi001;
assign w217 = pi053 & ~pi060;
assign w218 = w91 & w38;
assign w219 = w314 & w256;
assign w220 = ~pi031 & ~pi036;
assign w221 = ~pi062 & pi063;
assign w222 = ~w188 & ~pi025;
assign w223 = ~pi012 & pi037;
assign w224 = pi005 & w251;
assign w225 = ~pi014 & pi037;
assign w226 = ~pi037 & pi112;
assign w227 = ~pi095 & ~pi004;
assign w228 = (~pi029 & ~w85) | (~pi029 & w310) | (~w85 & w310);
assign w229 = w244 & w127;
assign w230 = pi039 & ~w20;
assign w231 = pi021 & ~pi018;
assign w232 = w73 & w298;
assign w233 = pi099 & ~w213;
assign w234 = pi038 & ~pi073;
assign w235 = pi058 & w265;
assign w236 = pi028 & w77;
assign w237 = w100 & ~w112;
assign w238 = (~w249 & ~w261) | (~w249 & w175) | (~w261 & w175);
assign w239 = w315 & w347;
assign w240 = ~w155 & ~w286;
assign w241 = ~pi039 & w20;
assign w242 = pi019 & ~w50;
assign w243 = pi099 & ~w37;
assign w244 = w328 & w168;
assign w245 = ~pi091 & w369;
assign w246 = ~pi035 & ~w91;
assign w247 = ~pi074 & ~w263;
assign w248 = ~pi069 & ~pi073;
assign w249 = ~pi017 & pi027;
assign w250 = pi061 & ~pi073;
assign w251 = (pi099 & ~w244) | (pi099 & w330) | (~w244 & w330);
assign w252 = w311 & w297;
assign w253 = ~w304 & ~w142;
assign w254 = ~w111 & ~w217;
assign w255 = pi068 & w293;
assign w256 = pi027 & pi060;
assign w257 = w232 & w188;
assign w258 = (~w80 & w46) | (~w80 & ~w144) | (w46 & ~w144);
assign w259 = ~pi058 & ~pi054;
assign w260 = pi073 & pi028;
assign w261 = ~pi091 & w32;
assign w262 = ~w168 & ~pi001;
assign w263 = ~pi083 & pi087;
assign w264 = ~w20 & w269;
assign w265 = pi026 & pi054;
assign w266 = ~w52 & ~w284;
assign w267 = ~pi037 & ~pi109;
assign w268 = ~w264 & w118;
assign w269 = pi039 & pi038;
assign w270 = ~w132 & w62;
assign w271 = ~pi026 & ~w232;
assign w272 = ~pi035 & w77;
assign w273 = w334 & ~w335;
assign w274 = ~pi073 & ~pi075;
assign w275 = (~pi043 & w264) | (~pi043 & w324) | (w264 & w324);
assign w276 = ~w274 & ~w354;
assign w277 = ~w291 & w79;
assign w278 = (~w50 & w238) | (~w50 & w242) | (w238 & w242);
assign w279 = pi060 & pi100;
assign w280 = pi028 & pi029;
assign w281 = pi062 & ~pi063;
assign w282 = ~w285 & w98;
assign w283 = (pi032 & ~w185) | (pi032 & w194) | (~w185 & w194);
assign w284 = ~pi011 & pi037;
assign w285 = ~w230 & ~w241;
assign w286 = w91 & w56;
assign w287 = ~pi037 & ~pi108;
assign w288 = ~pi062 & ~pi063;
assign w289 = ~w326 & w148;
assign w290 = ~pi004 & ~pi005;
assign w291 = ~pi069 & w48;
assign w292 = ~pi073 & w311;
assign w293 = ~pi073 & pi099;
assign w294 = ~w173 & ~pi042;
assign w295 = ~pi017 & ~pi019;
assign w296 = ~pi037 & ~pi105;
assign w297 = ~pi073 & pi039;
assign w298 = pi058 & pi054;
assign w299 = ~w261 & w332;
assign w300 = pi073 & ~w218;
assign w301 = ~w306 & w15;
assign w302 = pi065 & w63;
assign w303 = ~pi071 & pi100;
assign w304 = ~pi037 & ~pi106;
assign w305 = (~pi031 & ~w91) | (~pi031 & w86) | (~w91 & w86);
assign w306 = (~pi042 & w264) | (~pi042 & w294) | (w264 & w294);
assign w307 = ~w261 & ~w178;
assign w308 = pi095 & ~pi001;
assign w309 = pi097 & w198;
assign w310 = ~pi056 & ~pi029;
assign w311 = pi065 & pi099;
assign w312 = ~pi034 & w280;
assign w313 = pi056 & ~w288;
assign w314 = pi017 & ~pi019;
assign w315 = ~pi060 & pi073;
assign w316 = ~w110 & w1;
assign w317 = ~pi009 & pi037;
assign w318 = ~pi005 & ~w290;
assign w319 = pi099 & ~w365;
assign w320 = pi099 & ~w71;
assign w321 = pi019 & pi073;
assign w322 = ~w325 & w77;
assign w323 = pi092 & w198;
assign w324 = ~w190 & ~pi043;
assign w325 = pi035 & pi036;
assign w326 = (~pi036 & ~w91) | (~pi036 & w368) | (~w91 & w368);
assign w327 = ~w89 & ~w101;
assign w328 = pi073 & ~w288;
assign w329 = ~w147 & ~w154;
assign w330 = w49 & pi099;
assign w331 = pi099 & ~w95;
assign w332 = w146 & ~w321;
assign w333 = (w77 & w4) | (w77 & w236) | (w4 & w236);
assign w334 = pi099 & w212;
assign w335 = (~pi024 & ~w232) | (~pi024 & w123) | (~w232 & w123);
assign w336 = pi071 & ~w174;
assign w337 = pi018 & ~pi021;
assign w338 = ~w267 & ~w200;
assign w339 = w334 & ~w232;
assign w340 = pi004 & ~w251;
assign w341 = pi095 & w221;
assign w342 = pi060 & ~w164;
assign w343 = pi071 & ~w279;
assign w344 = ~w347 & ~w219;
assign w345 = pi065 & ~w184;
assign w346 = ~w282 & ~w252;
assign w347 = ~w6 & w151;
assign w348 = ~w246 & w143;
assign w349 = pi066 & w311;
assign w350 = ~w296 & ~w317;
assign w351 = pi000 & ~pi073;
assign w352 = ~w224 & ~w172;
assign w353 = (~w124 & w141) | (~w124 & w233) | (w141 & w233);
assign w354 = pi073 & ~pi074;
assign w355 = w244 & w11;
assign w356 = ~w275 & w358;
assign w357 = ~w42 & w26;
assign w358 = w311 & ~w183;
assign w359 = pi099 & ~w54;
assign w360 = ~w111 & w92;
assign w361 = ~w203 & w353;
assign w362 = pi067 & w293;
assign w363 = ~pi073 & ~pi041;
assign w364 = pi099 & ~w315;
assign w365 = (~w178 & ~w7) | (~w178 & w307) | (~w7 & w307);
assign w366 = ~w264 & w109;
assign w367 = ~pi071 & w174;
assign w368 = ~pi035 & ~pi036;
assign w369 = pi064 & pi077;
assign w370 = pi068 & pi073;
assign w371 = ~w64 & w333;
assign one = 1;
assign po000 = pi070;
assign po001 = pi055;
assign po002 = pi059;
assign po003 = pi061;
assign po004 = pi040;
assign po005 = pi044;
assign po006 = pi002;
assign po007 = ~w197;
assign po008 = pi047;
assign po009 = pi048;
assign po010 = pi049;
assign po011 = pi050;
assign po012 = pi046;
assign po013 = pi051;
assign po014 = pi045;
assign po015 = pi052;
assign po016 = pi084;
assign po017 = pi082;
assign po018 = one;
assign po019 = pi098;
assign po020 = ~w27;
assign po021 = w66;
assign po022 = w243;
assign po023 = w114;
assign po024 = w108;
assign po025 = ~w352;
assign po026 = w30;
assign po027 = ~w104;
assign po028 = w125;
assign po029 = w9;
assign po030 = w105;
assign po031 = w60;
assign po032 = w36;
assign po033 = w81;
assign po034 = w360;
assign po035 = w96;
assign po036 = w181;
assign po037 = w320;
assign po038 = ~w361;
assign po039 = w68;
assign po040 = w61;
assign po041 = w128;
assign po042 = ~w119;
assign po043 = w288;
assign po044 = w51;
assign po045 = w270;
assign po046 = w196;
assign po047 = w23;
assign po048 = w371;
assign po049 = w176;
assign po050 = w191;
assign po051 = w192;
assign po052 = w316;
assign po053 = w319;
assign po054 = w357;
assign po055 = w348;
assign po056 = w289;
assign po057 = w129;
assign po058 = w170;
assign po059 = ~w346;
assign po060 = w14;
assign po061 = w33;
assign po062 = w301;
assign po063 = w356;
assign po064 = w133;
assign po065 = ~w169;
assign po066 = pi056;
assign po067 = w130;
assign po068 = w93;
assign po069 = w329;
assign po070 = w331;
assign po071 = ~w163;
assign po072 = w84;
assign po073 = w76;
assign po074 = w359;
assign po075 = ~w277;
assign po076 = ~w28;
assign po077 = ~w34;
assign po078 = w366;
assign po079 = ~w106;
assign po080 = ~w149;
assign po081 = ~w102;
assign po082 = ~w69;
assign po083 = w208;
assign po084 = w214;
assign po085 = ~w74;
assign po086 = w120;
assign po087 = pi076;
assign po088 = w206;
assign po089 = w276;
assign po090 = pi080;
assign po091 = w237;
assign po092 = w16;
assign po093 = w31;
assign po094 = w337;
assign po095 = pi074;
assign po096 = pi089;
assign po097 = pi087;
assign po098 = pi093;
assign po099 = pi010;
assign po100 = pi014;
assign po101 = pi101;
assign po102 = pi012;
assign po103 = pi103;
assign po104 = pi015;
assign po105 = pi064;
assign po106 = pi009;
assign po107 = pi102;
assign po108 = pi011;
assign po109 = pi007;
assign po110 = pi013;
endmodule

// Benchmark "top" written by ABC on Tue Feb 13 00:53:45 2018

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110;
  wire n225, n226, n227, n228, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n306, n307, n308, n309, n310, n311, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n324, n325, n327, n328, n329,
    n330, n331, n332, n333, n334, n336, n337, n338, n339, n340, n341, n342,
    n343, n345, n346, n348, n349, n351, n352, n354, n355, n357, n358, n360,
    n361, n363, n364, n366, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n396, n397, n398, n399, n400,
    n401, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n414,
    n415, n416, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434, n436, n437, n438, n439, n440,
    n441, n443, n444, n445, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n468, n469, n470, n471, n472, n473, n474, n476, n477, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n505, n506, n507,
    n508, n509, n510, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n547, n548, n549, n550, n551, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, n571,
    n572, n573, n574, n576, n577, n578, n579, n580, n582, n583, n584, n585,
    n586, n587, n588, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n602, n603, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n615, n616, n617, n618, n619, n620, n621, n622, n624, n625, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n640,
    n641, n642, n643, n644, n646, n647, n648, n649, n650, n651, n654, n656,
    n657, n658, n660, n661, n662, n663, n664, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n677, n678, n679, n680, n681, n682, n683,
    n685, n686, n687, n689, n690, n692, n693, n694, n695, n696, n697, n699,
    n700, n701, n702, n703, n704, n706, n707, n708, n709, n711, n712, n713,
    n715, n717, n718, n719, n721, n724, n725, n726, n728, n729, n730, n731,
    n733, n734, n735, n736, n738, n739, n740, n742, n743, n745, n746, n748,
    n749, n750, n751, n753, n755, n756, n757, n758, n759, n761, n762, n764;
  inv1 g000(.a(pi003), .O(n225));
  inv1 g001(.a(pi006), .O(n226));
  inv1 g002(.a(pi008), .O(n227));
  nor3 g003(.a(n227), .b(n226), .c(n225), .O(n228));
  inv1 g004(.a(n228), .O(po007));
  inv1 g005(.a(pi005), .O(n231));
  inv1 g006(.a(pi062), .O(n232));
  nor2 g007(.a(pi095), .b(pi004), .O(n233));
  nor3 g008(.a(n233), .b(pi063), .c(n232), .O(n234));
  nor2 g009(.a(n234), .b(pi004), .O(n235));
  nor2 g010(.a(pi063), .b(n232), .O(n236));
  inv1 g011(.a(n233), .O(n237));
  nor2 g012(.a(n237), .b(n236), .O(n238));
  nor3 g013(.a(n238), .b(n235), .c(n231), .O(n239));
  inv1 g014(.a(n239), .O(n240));
  inv1 g015(.a(pi001), .O(n241));
  inv1 g016(.a(n236), .O(n242));
  inv1 g017(.a(pi073), .O(n243));
  nor2 g018(.a(pi063), .b(pi062), .O(po043));
  nor2 g019(.a(po043), .b(n243), .O(n245));
  inv1 g020(.a(n245), .O(n246));
  nor2 g021(.a(pi016), .b(pi002), .O(n247));
  inv1 g022(.a(n247), .O(n248));
  nor2 g023(.a(n248), .b(n246), .O(n249));
  inv1 g024(.a(n249), .O(n250));
  nor3 g025(.a(n250), .b(n242), .c(n241), .O(n251));
  inv1 g026(.a(n251), .O(n252));
  nor2 g027(.a(n252), .b(n240), .O(n253));
  inv1 g028(.a(pi000), .O(n254));
  nor2 g029(.a(pi073), .b(n254), .O(n255));
  inv1 g030(.a(pi002), .O(n256));
  nor2 g031(.a(n243), .b(n256), .O(n257));
  nor3 g032(.a(n257), .b(n255), .c(n253), .O(n258));
  inv1 g033(.a(n258), .O(po020));
  nor2 g034(.a(n247), .b(pi001), .O(n260));
  nor2 g035(.a(n260), .b(n246), .O(n261));
  nor2 g036(.a(n261), .b(pi001), .O(n262));
  inv1 g037(.a(n260), .O(n263));
  nor2 g038(.a(n263), .b(n245), .O(n264));
  inv1 g039(.a(pi099), .O(n265));
  inv1 g040(.a(pi095), .O(n266));
  nor3 g041(.a(n242), .b(n266), .c(pi001), .O(n267));
  inv1 g042(.a(n267), .O(n268));
  nor3 g043(.a(n268), .b(n249), .c(n265), .O(n269));
  nor2 g044(.a(n268), .b(n265), .O(n270));
  nor2 g045(.a(n270), .b(n250), .O(n271));
  nor2 g046(.a(n271), .b(n265), .O(n272));
  nor2 g047(.a(n272), .b(n269), .O(n273));
  nor3 g048(.a(n273), .b(n264), .c(n262), .O(po021));
  nor3 g049(.a(po043), .b(pi022), .c(n256), .O(n275));
  inv1 g050(.a(po043), .O(n276));
  nor2 g051(.a(pi022), .b(n256), .O(n277));
  nor2 g052(.a(n277), .b(n276), .O(n278));
  nor2 g053(.a(n278), .b(n256), .O(n279));
  nor2 g054(.a(n279), .b(n275), .O(n280));
  nor3 g055(.a(n279), .b(n275), .c(pi095), .O(n281));
  nor2 g056(.a(n281), .b(n280), .O(n282));
  inv1 g057(.a(n280), .O(n283));
  nor2 g058(.a(n281), .b(n240), .O(n284));
  nor2 g059(.a(n284), .b(n283), .O(n285));
  inv1 g060(.a(n281), .O(n286));
  nor2 g061(.a(n286), .b(n239), .O(n287));
  nor2 g062(.a(n287), .b(n285), .O(n288));
  nor2 g063(.a(n288), .b(n282), .O(n289));
  inv1 g064(.a(n282), .O(n290));
  nor3 g065(.a(n287), .b(n285), .c(n290), .O(n291));
  nor2 g066(.a(n291), .b(n251), .O(n292));
  nor3 g067(.a(n292), .b(n289), .c(n265), .O(po022));
  inv1 g068(.a(pi063), .O(n294));
  nor2 g069(.a(n294), .b(pi062), .O(n295));
  inv1 g070(.a(n295), .O(n296));
  nor3 g071(.a(n296), .b(n266), .c(n241), .O(n297));
  nor2 g072(.a(n297), .b(n239), .O(n298));
  nor2 g073(.a(n298), .b(n241), .O(n299));
  inv1 g074(.a(n297), .O(n300));
  nor2 g075(.a(n300), .b(n240), .O(n301));
  nor3 g076(.a(pi005), .b(pi004), .c(pi001), .O(n302));
  nor3 g077(.a(n302), .b(n267), .c(n250), .O(n303));
  inv1 g078(.a(n303), .O(n304));
  nor3 g079(.a(n304), .b(n301), .c(n299), .O(po023));
  nor4 g080(.a(n296), .b(n265), .c(n266), .d(n241), .O(n306));
  inv1 g081(.a(n306), .O(n307));
  nor2 g082(.a(n307), .b(n250), .O(n308));
  nor2 g083(.a(n308), .b(pi004), .O(n309));
  inv1 g084(.a(pi004), .O(n310));
  nor3 g085(.a(n272), .b(n269), .c(n310), .O(n311));
  nor2 g086(.a(n311), .b(n309), .O(po024));
  nor2 g087(.a(n273), .b(n231), .O(n313));
  inv1 g088(.a(n308), .O(n314));
  nor4 g089(.a(n237), .b(n236), .c(pi005), .d(n310), .O(n315));
  nor2 g090(.a(pi005), .b(pi004), .O(n316));
  nor2 g091(.a(pi005), .b(n310), .O(n317));
  nor3 g092(.a(n317), .b(n238), .c(n235), .O(n318));
  nor2 g093(.a(n318), .b(n316), .O(n319));
  nor2 g094(.a(n319), .b(n315), .O(n320));
  nor2 g095(.a(n320), .b(n314), .O(n321));
  nor2 g096(.a(n321), .b(n313), .O(n322));
  inv1 g097(.a(n322), .O(po025));
  inv1 g098(.a(pi023), .O(n324));
  nor2 g099(.a(pi036), .b(pi031), .O(n325));
  nor4 g100(.a(n325), .b(n276), .c(n324), .d(n256), .O(po026));
  inv1 g101(.a(pi104), .O(n327));
  nor4 g102(.a(n327), .b(pi027), .c(pi019), .d(pi017), .O(n328));
  inv1 g103(.a(pi112), .O(n329));
  nor2 g104(.a(n329), .b(pi037), .O(n330));
  inv1 g105(.a(pi007), .O(n331));
  inv1 g106(.a(pi037), .O(n332));
  nor2 g107(.a(n332), .b(n331), .O(n333));
  nor3 g108(.a(n333), .b(n330), .c(n328), .O(n334));
  inv1 g109(.a(n334), .O(po027));
  inv1 g110(.a(n257), .O(n336));
  inv1 g111(.a(pi028), .O(n337));
  inv1 g112(.a(pi029), .O(n338));
  nor2 g113(.a(n338), .b(n337), .O(n339));
  inv1 g114(.a(n339), .O(n340));
  inv1 g115(.a(pi056), .O(n341));
  nor2 g116(.a(po043), .b(n341), .O(n342));
  inv1 g117(.a(n342), .O(n343));
  nor4 g118(.a(n343), .b(n340), .c(n336), .d(pi034), .O(po028));
  nor2 g119(.a(pi105), .b(pi037), .O(n345));
  nor2 g120(.a(n332), .b(pi009), .O(n346));
  nor3 g121(.a(n346), .b(n345), .c(n328), .O(po029));
  nor2 g122(.a(pi106), .b(pi037), .O(n348));
  nor2 g123(.a(n332), .b(pi010), .O(n349));
  nor3 g124(.a(n349), .b(n348), .c(n328), .O(po030));
  nor2 g125(.a(pi107), .b(pi037), .O(n351));
  nor2 g126(.a(n332), .b(pi011), .O(n352));
  nor3 g127(.a(n352), .b(n351), .c(n328), .O(po031));
  nor2 g128(.a(pi108), .b(pi037), .O(n354));
  nor2 g129(.a(n332), .b(pi012), .O(n355));
  nor3 g130(.a(n355), .b(n354), .c(n328), .O(po032));
  nor2 g131(.a(pi109), .b(pi037), .O(n357));
  nor2 g132(.a(n332), .b(pi013), .O(n358));
  nor3 g133(.a(n358), .b(n357), .c(n328), .O(po033));
  nor2 g134(.a(pi110), .b(pi037), .O(n360));
  nor2 g135(.a(n332), .b(pi014), .O(n361));
  nor3 g136(.a(n361), .b(n360), .c(n328), .O(po034));
  nor2 g137(.a(pi111), .b(pi037), .O(n363));
  nor2 g138(.a(n332), .b(pi015), .O(n364));
  nor3 g139(.a(n364), .b(n363), .c(n328), .O(po035));
  nor2 g140(.a(pi073), .b(pi016), .O(n366));
  nor2 g141(.a(n366), .b(n245), .O(po036));
  inv1 g142(.a(pi064), .O(n368));
  nor3 g143(.a(pi091), .b(n368), .c(pi019), .O(n369));
  inv1 g144(.a(n369), .O(n370));
  inv1 g145(.a(pi077), .O(n371));
  nor3 g146(.a(pi091), .b(n371), .c(n368), .O(n372));
  inv1 g147(.a(pi027), .O(n373));
  nor2 g148(.a(n373), .b(pi017), .O(n374));
  inv1 g149(.a(n374), .O(n375));
  nor2 g150(.a(n375), .b(n372), .O(n376));
  inv1 g151(.a(n376), .O(n377));
  nor2 g152(.a(n377), .b(n370), .O(n378));
  inv1 g153(.a(pi017), .O(n379));
  nor4 g154(.a(pi060), .b(n373), .c(pi019), .d(n379), .O(n380));
  nor2 g155(.a(n380), .b(n328), .O(n381));
  inv1 g156(.a(n381), .O(n382));
  inv1 g157(.a(pi019), .O(n383));
  nor2 g158(.a(n243), .b(n383), .O(n384));
  nor2 g159(.a(pi027), .b(n379), .O(n385));
  inv1 g160(.a(n385), .O(n386));
  nor3 g161(.a(n386), .b(n384), .c(n369), .O(n387));
  nor2 g162(.a(n243), .b(pi060), .O(n388));
  inv1 g163(.a(n388), .O(n389));
  nor2 g164(.a(n243), .b(n379), .O(n390));
  nor3 g165(.a(n390), .b(pi027), .c(n383), .O(n391));
  inv1 g166(.a(n391), .O(n392));
  nor2 g167(.a(n392), .b(n389), .O(n393));
  nor4 g168(.a(n393), .b(n387), .c(n382), .d(n378), .O(n394));
  nor2 g169(.a(n394), .b(n265), .O(po037));
  inv1 g170(.a(pi081), .O(n396));
  nor2 g171(.a(n396), .b(pi074), .O(n397));
  inv1 g172(.a(pi074), .O(n398));
  nor2 g173(.a(pi081), .b(n398), .O(n399));
  nor2 g174(.a(n399), .b(n397), .O(n400));
  inv1 g175(.a(pi018), .O(n401));
  nor2 g176(.a(pi021), .b(n401), .O(po094));
  inv1 g177(.a(po094), .O(n403));
  nor3 g178(.a(n403), .b(n400), .c(n266), .O(n404));
  nor2 g179(.a(pi095), .b(pi018), .O(n405));
  nor3 g180(.a(n405), .b(n265), .c(n401), .O(n406));
  nor2 g181(.a(n265), .b(n401), .O(n407));
  nor2 g182(.a(n405), .b(n265), .O(n408));
  nor2 g183(.a(n408), .b(n407), .O(n409));
  nor2 g184(.a(n409), .b(n400), .O(n410));
  nor2 g185(.a(n410), .b(n406), .O(n411));
  nor2 g186(.a(n411), .b(n404), .O(n412));
  inv1 g187(.a(n412), .O(po038));
  inv1 g188(.a(pi060), .O(n414));
  nor4 g189(.a(n414), .b(n373), .c(pi019), .d(n379), .O(n415));
  nor2 g190(.a(n415), .b(n391), .O(n416));
  nor2 g191(.a(n416), .b(n265), .O(po039));
  inv1 g192(.a(pi020), .O(n418));
  inv1 g193(.a(pi034), .O(n419));
  nor2 g194(.a(n243), .b(n419), .O(n420));
  inv1 g195(.a(n420), .O(n421));
  nor2 g196(.a(n421), .b(n339), .O(n422));
  nor2 g197(.a(n420), .b(n340), .O(n423));
  nor2 g198(.a(n423), .b(n243), .O(n424));
  nor2 g199(.a(n424), .b(n422), .O(n425));
  inv1 g200(.a(n425), .O(n426));
  nor2 g201(.a(n426), .b(n418), .O(n427));
  inv1 g202(.a(pi031), .O(n428));
  inv1 g203(.a(pi035), .O(n429));
  inv1 g204(.a(pi036), .O(n430));
  nor2 g205(.a(n430), .b(n429), .O(n431));
  inv1 g206(.a(n431), .O(n432));
  nor3 g207(.a(n432), .b(n425), .c(n428), .O(n433));
  nor2 g208(.a(n433), .b(n427), .O(n434));
  nor2 g209(.a(n434), .b(n265), .O(po040));
  inv1 g210(.a(pi021), .O(n436));
  nor2 g211(.a(n436), .b(pi018), .O(n437));
  inv1 g212(.a(n437), .O(n438));
  nor3 g213(.a(n438), .b(n399), .c(n397), .O(n439));
  nor3 g214(.a(pi095), .b(n436), .c(pi018), .O(n440));
  nor3 g215(.a(n440), .b(n439), .c(po094), .O(n441));
  nor2 g216(.a(n441), .b(n265), .O(po041));
  inv1 g217(.a(pi022), .O(n443));
  nor2 g218(.a(pi073), .b(n443), .O(n444));
  nor2 g219(.a(n444), .b(pi044), .O(n445));
  inv1 g220(.a(n445), .O(po042));
  nor2 g221(.a(n243), .b(pi070), .O(n447));
  inv1 g222(.a(n447), .O(n448));
  inv1 g223(.a(pi054), .O(n449));
  inv1 g224(.a(pi058), .O(n450));
  nor2 g225(.a(n450), .b(n449), .O(n451));
  inv1 g226(.a(n451), .O(n452));
  nor2 g227(.a(n452), .b(n448), .O(n453));
  inv1 g228(.a(n453), .O(n454));
  inv1 g229(.a(pi024), .O(n455));
  inv1 g230(.a(pi026), .O(n456));
  nor2 g231(.a(n456), .b(n455), .O(n457));
  inv1 g232(.a(n457), .O(n458));
  nor2 g233(.a(n458), .b(n454), .O(n459));
  nor2 g234(.a(pi026), .b(pi024), .O(n460));
  nor2 g235(.a(n460), .b(n454), .O(n461));
  nor2 g236(.a(n461), .b(pi024), .O(n462));
  inv1 g237(.a(n460), .O(n463));
  nor2 g238(.a(n463), .b(n453), .O(n464));
  nor3 g239(.a(n265), .b(pi084), .c(pi082), .O(n465));
  inv1 g240(.a(n465), .O(n466));
  nor4 g241(.a(n466), .b(n464), .c(n462), .d(n459), .O(po044));
  inv1 g242(.a(pi025), .O(n468));
  nor3 g243(.a(n458), .b(n454), .c(n468), .O(n469));
  nor2 g244(.a(n457), .b(pi025), .O(n470));
  nor2 g245(.a(n470), .b(n454), .O(n471));
  nor2 g246(.a(n471), .b(pi025), .O(n472));
  inv1 g247(.a(n470), .O(n473));
  nor2 g248(.a(n473), .b(n453), .O(n474));
  nor4 g249(.a(n474), .b(n472), .c(n469), .d(n466), .O(po045));
  nor2 g250(.a(n453), .b(pi026), .O(n476));
  nor2 g251(.a(n454), .b(n456), .O(n477));
  nor3 g252(.a(n477), .b(n476), .c(n466), .O(po046));
  nor2 g253(.a(n385), .b(n374), .O(n479));
  nor2 g254(.a(n479), .b(n370), .O(n480));
  nor2 g255(.a(n480), .b(n374), .O(n481));
  nor3 g256(.a(n385), .b(n374), .c(n369), .O(n482));
  nor2 g257(.a(n482), .b(n481), .O(n483));
  nor2 g258(.a(n380), .b(n383), .O(n484));
  inv1 g259(.a(n484), .O(n485));
  nor2 g260(.a(n485), .b(n483), .O(n486));
  inv1 g261(.a(n483), .O(n487));
  nor2 g262(.a(n484), .b(n487), .O(n488));
  nor2 g263(.a(n488), .b(n380), .O(n489));
  nor3 g264(.a(n489), .b(n486), .c(n265), .O(po047));
  nor2 g265(.a(n419), .b(n338), .O(n491));
  nor3 g266(.a(n491), .b(n425), .c(n341), .O(n492));
  nor3 g267(.a(n492), .b(n243), .c(n337), .O(n493));
  nor2 g268(.a(n265), .b(n254), .O(n494));
  inv1 g269(.a(n494), .O(n495));
  nor4 g270(.a(n243), .b(n341), .c(n419), .d(n338), .O(n496));
  nor2 g271(.a(n495), .b(n337), .O(n497));
  nor2 g272(.a(n497), .b(n496), .O(n498));
  nor2 g273(.a(n498), .b(n495), .O(n499));
  inv1 g274(.a(n496), .O(n500));
  inv1 g275(.a(n497), .O(n501));
  nor2 g276(.a(n501), .b(n500), .O(n502));
  nor2 g277(.a(n502), .b(n499), .O(n503));
  nor2 g278(.a(n503), .b(n493), .O(po048));
  nor2 g279(.a(n492), .b(n243), .O(n505));
  nor2 g280(.a(pi056), .b(pi029), .O(n506));
  nor2 g281(.a(n506), .b(n421), .O(n507));
  nor2 g282(.a(n507), .b(pi029), .O(n508));
  inv1 g283(.a(n506), .O(n509));
  nor2 g284(.a(n509), .b(n420), .O(n510));
  nor4 g285(.a(n510), .b(n508), .c(n505), .d(n495), .O(po049));
  inv1 g286(.a(pi065), .O(n512));
  inv1 g287(.a(pi041), .O(n513));
  nor2 g288(.a(pi042), .b(n513), .O(n514));
  inv1 g289(.a(n514), .O(n515));
  nor2 g290(.a(n515), .b(pi085), .O(n516));
  inv1 g291(.a(pi042), .O(n517));
  inv1 g292(.a(pi094), .O(n518));
  nor3 g293(.a(n518), .b(n517), .c(pi041), .O(n519));
  inv1 g294(.a(pi092), .O(n520));
  nor3 g295(.a(n520), .b(pi042), .c(pi041), .O(n521));
  nor2 g296(.a(n517), .b(n513), .O(n522));
  inv1 g297(.a(n522), .O(n523));
  inv1 g298(.a(pi088), .O(n524));
  nor2 g299(.a(n524), .b(pi032), .O(n525));
  nor2 g300(.a(n525), .b(n523), .O(n526));
  nor2 g301(.a(n526), .b(pi032), .O(n527));
  inv1 g302(.a(n525), .O(n528));
  nor2 g303(.a(n528), .b(n522), .O(n529));
  nor2 g304(.a(n529), .b(n527), .O(n530));
  nor4 g305(.a(n530), .b(n521), .c(n519), .d(n516), .O(n531));
  inv1 g306(.a(pi096), .O(n532));
  nor2 g307(.a(n523), .b(n532), .O(n533));
  nor3 g308(.a(pi090), .b(n517), .c(pi041), .O(n534));
  inv1 g309(.a(pi097), .O(n535));
  nor3 g310(.a(n535), .b(pi042), .c(pi041), .O(n536));
  inv1 g311(.a(pi032), .O(n537));
  inv1 g312(.a(pi086), .O(n538));
  nor2 g313(.a(n538), .b(n537), .O(n539));
  inv1 g314(.a(n539), .O(n540));
  nor2 g315(.a(n540), .b(n514), .O(n541));
  nor2 g316(.a(n539), .b(n515), .O(n542));
  nor2 g317(.a(n542), .b(n537), .O(n543));
  nor2 g318(.a(n543), .b(n541), .O(n544));
  nor4 g319(.a(n544), .b(n536), .c(n534), .d(n533), .O(n545));
  nor3 g320(.a(n545), .b(n531), .c(n512), .O(po050));
  nor2 g321(.a(n431), .b(pi031), .O(n547));
  nor2 g322(.a(n547), .b(n425), .O(n548));
  nor2 g323(.a(n548), .b(pi031), .O(n549));
  inv1 g324(.a(n547), .O(n550));
  nor2 g325(.a(n550), .b(n426), .O(n551));
  nor4 g326(.a(n551), .b(n549), .c(n495), .d(n433), .O(po051));
  inv1 g327(.a(pi038), .O(n553));
  inv1 g328(.a(pi039), .O(n554));
  nor3 g329(.a(pi043), .b(n554), .c(n553), .O(n555));
  nor3 g330(.a(n555), .b(n523), .c(n243), .O(n556));
  inv1 g331(.a(n556), .O(n557));
  nor2 g332(.a(n557), .b(n537), .O(n558));
  nor2 g333(.a(n265), .b(n512), .O(n559));
  inv1 g334(.a(n559), .O(n560));
  nor2 g335(.a(n560), .b(n537), .O(n561));
  nor2 g336(.a(n561), .b(n556), .O(n562));
  nor2 g337(.a(n562), .b(n560), .O(n563));
  inv1 g338(.a(n561), .O(n564));
  nor2 g339(.a(n564), .b(n557), .O(n565));
  nor2 g340(.a(n565), .b(n563), .O(n566));
  nor2 g341(.a(n566), .b(n558), .O(po052));
  inv1 g342(.a(pi033), .O(n568));
  nor2 g343(.a(pi068), .b(n568), .O(n569));
  nor2 g344(.a(n569), .b(n369), .O(n570));
  nor2 g345(.a(n570), .b(n377), .O(n571));
  nor2 g346(.a(n571), .b(n569), .O(n572));
  inv1 g347(.a(n570), .O(n573));
  nor2 g348(.a(n573), .b(n376), .O(n574));
  nor3 g349(.a(n574), .b(n572), .c(n265), .O(po053));
  nor2 g350(.a(pi056), .b(pi034), .O(n576));
  nor2 g351(.a(n576), .b(n425), .O(n577));
  nor2 g352(.a(n577), .b(pi034), .O(n578));
  inv1 g353(.a(n576), .O(n579));
  nor2 g354(.a(n579), .b(n426), .O(n580));
  nor4 g355(.a(n580), .b(n578), .c(n495), .d(n420), .O(po054));
  nor2 g356(.a(n426), .b(pi035), .O(n582));
  nor2 g357(.a(n495), .b(pi035), .O(n583));
  inv1 g358(.a(n583), .O(n584));
  nor2 g359(.a(n584), .b(n426), .O(n585));
  nor2 g360(.a(n583), .b(n425), .O(n586));
  nor2 g361(.a(n586), .b(n495), .O(n587));
  nor2 g362(.a(n587), .b(n585), .O(n588));
  nor2 g363(.a(n588), .b(n582), .O(po055));
  nor2 g364(.a(pi036), .b(pi035), .O(n590));
  nor2 g365(.a(n590), .b(n425), .O(n591));
  nor2 g366(.a(n591), .b(pi036), .O(n592));
  inv1 g367(.a(n590), .O(n593));
  nor2 g368(.a(n593), .b(n426), .O(n594));
  nor2 g369(.a(n495), .b(n431), .O(n595));
  inv1 g370(.a(n595), .O(n596));
  nor2 g371(.a(n596), .b(n426), .O(n597));
  nor2 g372(.a(n595), .b(n425), .O(n598));
  nor2 g373(.a(n598), .b(n495), .O(n599));
  nor2 g374(.a(n599), .b(n597), .O(n600));
  nor3 g375(.a(n600), .b(n594), .c(n592), .O(po056));
  nor2 g376(.a(n487), .b(n376), .O(n602));
  inv1 g377(.a(n602), .O(n603));
  nor3 g378(.a(n603), .b(n368), .c(pi019), .O(po057));
  nor2 g379(.a(pi073), .b(n553), .O(n605));
  inv1 g380(.a(pi043), .O(n606));
  nor2 g381(.a(n606), .b(n553), .O(n607));
  inv1 g382(.a(pi030), .O(n608));
  nor2 g383(.a(n243), .b(n608), .O(n609));
  inv1 g384(.a(n609), .O(n610));
  nor3 g385(.a(n610), .b(n555), .c(n607), .O(n611));
  nor2 g386(.a(n611), .b(n605), .O(n612));
  nor2 g387(.a(pi043), .b(pi038), .O(n613));
  nor3 g388(.a(n613), .b(n612), .c(n560), .O(po058));
  nor2 g389(.a(n607), .b(n554), .O(n615));
  nor3 g390(.a(n606), .b(pi039), .c(n553), .O(n616));
  nor2 g391(.a(n616), .b(n615), .O(n617));
  nor3 g392(.a(n610), .b(n560), .c(n555), .O(n618));
  inv1 g393(.a(n618), .O(n619));
  nor2 g394(.a(n619), .b(n617), .O(n620));
  nor3 g395(.a(n560), .b(pi073), .c(n554), .O(n621));
  nor2 g396(.a(n621), .b(n620), .O(n622));
  inv1 g397(.a(n622), .O(po059));
  nor2 g398(.a(n327), .b(n265), .O(n624));
  inv1 g399(.a(n624), .O(n625));
  nor2 g400(.a(n625), .b(n603), .O(po060));
  inv1 g401(.a(n555), .O(n627));
  nor2 g402(.a(pi073), .b(pi041), .O(n628));
  inv1 g403(.a(n628), .O(n629));
  nor2 g404(.a(n629), .b(n627), .O(n630));
  nor2 g405(.a(n628), .b(n555), .O(n631));
  nor2 g406(.a(n631), .b(pi041), .O(n632));
  nor2 g407(.a(n243), .b(n513), .O(n633));
  nor2 g408(.a(n633), .b(n560), .O(n634));
  nor2 g409(.a(n634), .b(n555), .O(n635));
  nor2 g410(.a(n635), .b(n560), .O(n636));
  nor3 g411(.a(n633), .b(n560), .c(n627), .O(n637));
  nor2 g412(.a(n637), .b(n636), .O(n638));
  nor3 g413(.a(n638), .b(n632), .c(n630), .O(po061));
  nor2 g414(.a(n633), .b(pi042), .O(n640));
  inv1 g415(.a(n640), .O(n641));
  nor2 g416(.a(n641), .b(n627), .O(n642));
  nor2 g417(.a(n640), .b(n555), .O(n643));
  nor2 g418(.a(n643), .b(pi042), .O(n644));
  nor4 g419(.a(n644), .b(n642), .c(n560), .d(n556), .O(po062));
  nor2 g420(.a(n609), .b(pi043), .O(n646));
  inv1 g421(.a(n646), .O(n647));
  nor2 g422(.a(n647), .b(n627), .O(n648));
  nor2 g423(.a(n646), .b(n555), .O(n649));
  nor2 g424(.a(n649), .b(pi043), .O(n650));
  nor2 g425(.a(n243), .b(n606), .O(n651));
  nor4 g426(.a(n651), .b(n650), .c(n648), .d(n560), .O(po063));
  nor2 g427(.a(n425), .b(n418), .O(po064));
  nor2 g428(.a(n425), .b(n254), .O(n654));
  inv1 g429(.a(n654), .O(po065));
  inv1 g430(.a(pi053), .O(n656));
  nor2 g431(.a(pi060), .b(n656), .O(n657));
  nor2 g432(.a(n657), .b(n328), .O(n658));
  nor2 g433(.a(n658), .b(n265), .O(po067));
  nor2 g434(.a(pi058), .b(pi054), .O(n660));
  nor2 g435(.a(n660), .b(n448), .O(n661));
  nor2 g436(.a(n661), .b(pi054), .O(n662));
  inv1 g437(.a(n660), .O(n663));
  nor2 g438(.a(n663), .b(n447), .O(n664));
  nor4 g439(.a(n664), .b(n662), .c(n466), .d(n453), .O(po068));
  nor2 g440(.a(n265), .b(pi073), .O(n666));
  inv1 g441(.a(n666), .O(n667));
  nor2 g442(.a(n667), .b(pi055), .O(n668));
  inv1 g443(.a(pi071), .O(n669));
  inv1 g444(.a(pi100), .O(n670));
  nor2 g445(.a(n670), .b(n414), .O(n671));
  nor2 g446(.a(n671), .b(n669), .O(n672));
  nor2 g447(.a(n265), .b(n243), .O(n673));
  inv1 g448(.a(n673), .O(n674));
  nor2 g449(.a(n674), .b(n672), .O(n675));
  nor2 g450(.a(n675), .b(n668), .O(po069));
  inv1 g451(.a(pi075), .O(n677));
  nor2 g452(.a(n677), .b(n398), .O(n678));
  nor2 g453(.a(pi075), .b(pi074), .O(n679));
  nor2 g454(.a(n679), .b(n678), .O(n680));
  nor2 g455(.a(n680), .b(n243), .O(n681));
  nor2 g456(.a(pi073), .b(n341), .O(n682));
  nor3 g457(.a(n682), .b(n681), .c(n256), .O(n683));
  nor2 g458(.a(n683), .b(n265), .O(po070));
  inv1 g459(.a(pi057), .O(n685));
  nor2 g460(.a(n667), .b(n685), .O(n686));
  nor2 g461(.a(n686), .b(n618), .O(n687));
  inv1 g462(.a(n687), .O(po071));
  nor2 g463(.a(n447), .b(pi058), .O(n689));
  nor2 g464(.a(n448), .b(n450), .O(n690));
  nor3 g465(.a(n690), .b(n689), .c(n466), .O(po072));
  nor2 g466(.a(n670), .b(pi071), .O(n692));
  nor2 g467(.a(n692), .b(n389), .O(n693));
  nor2 g468(.a(n674), .b(n671), .O(n694));
  inv1 g469(.a(pi059), .O(n695));
  nor2 g470(.a(n667), .b(n695), .O(n696));
  nor2 g471(.a(n696), .b(n694), .O(n697));
  nor2 g472(.a(n697), .b(n693), .O(po073));
  inv1 g473(.a(pi072), .O(n699));
  nor2 g474(.a(n243), .b(n699), .O(n700));
  nor2 g475(.a(n700), .b(n414), .O(n701));
  inv1 g476(.a(pi068), .O(n702));
  nor2 g477(.a(n243), .b(n702), .O(n703));
  nor2 g478(.a(n703), .b(n701), .O(n704));
  nor2 g479(.a(n704), .b(n265), .O(po074));
  nor3 g480(.a(n243), .b(pi069), .c(pi066), .O(n706));
  inv1 g481(.a(pi061), .O(n707));
  nor2 g482(.a(pi073), .b(n707), .O(n708));
  nor3 g483(.a(n708), .b(n706), .c(n265), .O(n709));
  inv1 g484(.a(n709), .O(po075));
  inv1 g485(.a(pi078), .O(n711));
  inv1 g486(.a(pi082), .O(n712));
  inv1 g487(.a(pi089), .O(n713));
  nor2 g488(.a(n713), .b(n712), .O(po092));
  nor2 g489(.a(po092), .b(n711), .O(n715));
  inv1 g490(.a(n715), .O(po076));
  inv1 g491(.a(pi079), .O(n717));
  inv1 g492(.a(pi084), .O(n718));
  inv1 g493(.a(pi093), .O(n719));
  nor2 g494(.a(n719), .b(n718), .O(po093));
  nor2 g495(.a(po093), .b(n717), .O(n721));
  inv1 g496(.a(n721), .O(po077));
  nor3 g497(.a(n555), .b(n523), .c(n537), .O(po078));
  nor2 g498(.a(n560), .b(pi073), .O(n724));
  nor2 g499(.a(n674), .b(n656), .O(n725));
  nor2 g500(.a(n725), .b(n724), .O(n726));
  inv1 g501(.a(n726), .O(po079));
  inv1 g502(.a(pi066), .O(n728));
  nor2 g503(.a(n667), .b(n728), .O(n729));
  nor2 g504(.a(n674), .b(n512), .O(n730));
  nor2 g505(.a(n730), .b(n729), .O(n731));
  inv1 g506(.a(n731), .O(po080));
  nor2 g507(.a(n674), .b(n568), .O(n733));
  inv1 g508(.a(pi067), .O(n734));
  nor2 g509(.a(n667), .b(n734), .O(n735));
  nor2 g510(.a(n735), .b(n733), .O(n736));
  inv1 g511(.a(n736), .O(po081));
  nor2 g512(.a(n674), .b(n734), .O(n738));
  nor2 g513(.a(n667), .b(n702), .O(n739));
  nor2 g514(.a(n739), .b(n738), .O(n740));
  inv1 g515(.a(n740), .O(po082));
  nor2 g516(.a(n243), .b(pi066), .O(n742));
  nor2 g517(.a(pi073), .b(pi069), .O(n743));
  nor3 g518(.a(n743), .b(n742), .c(n265), .O(po083));
  nor3 g519(.a(n450), .b(n449), .c(n456), .O(n745));
  inv1 g520(.a(n745), .O(n746));
  nor3 g521(.a(n746), .b(n468), .c(n455), .O(po084));
  nor3 g522(.a(n243), .b(pi071), .c(pi057), .O(n748));
  nor2 g523(.a(n243), .b(pi057), .O(n749));
  nor2 g524(.a(n749), .b(n669), .O(n750));
  nor4 g525(.a(n750), .b(n748), .c(n560), .d(n728), .O(n751));
  inv1 g526(.a(n751), .O(po085));
  nor2 g527(.a(pi073), .b(pi072), .O(n753));
  nor3 g528(.a(n753), .b(n388), .c(n265), .O(po086));
  inv1 g529(.a(pi083), .O(n755));
  nor2 g530(.a(pi087), .b(n755), .O(n756));
  inv1 g531(.a(pi087), .O(n757));
  nor2 g532(.a(n757), .b(pi083), .O(n758));
  nor2 g533(.a(n758), .b(pi074), .O(n759));
  nor2 g534(.a(n759), .b(n756), .O(po088));
  nor2 g535(.a(pi075), .b(pi073), .O(n761));
  nor2 g536(.a(pi074), .b(n243), .O(n762));
  nor2 g537(.a(n762), .b(n761), .O(po089));
  nor2 g538(.a(pi077), .b(n656), .O(n764));
  nor2 g539(.a(n764), .b(n625), .O(po091));
  one  g540(.O(po018));
  buf  g541(.a(pi070), .O(po000));
  buf  g542(.a(pi055), .O(po001));
  buf  g543(.a(pi059), .O(po002));
  buf  g544(.a(pi061), .O(po003));
  buf  g545(.a(pi040), .O(po004));
  buf  g546(.a(pi044), .O(po005));
  buf  g547(.a(pi002), .O(po006));
  buf  g548(.a(pi047), .O(po008));
  buf  g549(.a(pi048), .O(po009));
  buf  g550(.a(pi049), .O(po010));
  buf  g551(.a(pi050), .O(po011));
  buf  g552(.a(pi046), .O(po012));
  buf  g553(.a(pi051), .O(po013));
  buf  g554(.a(pi045), .O(po014));
  buf  g555(.a(pi052), .O(po015));
  buf  g556(.a(pi084), .O(po016));
  buf  g557(.a(pi082), .O(po017));
  buf  g558(.a(pi098), .O(po019));
  buf  g559(.a(pi056), .O(po066));
  buf  g560(.a(pi076), .O(po087));
  buf  g561(.a(pi080), .O(po090));
  buf  g562(.a(pi074), .O(po095));
  buf  g563(.a(pi089), .O(po096));
  buf  g564(.a(pi087), .O(po097));
  buf  g565(.a(pi093), .O(po098));
  buf  g566(.a(pi010), .O(po099));
  buf  g567(.a(pi014), .O(po100));
  buf  g568(.a(pi101), .O(po101));
  buf  g569(.a(pi012), .O(po102));
  buf  g570(.a(pi103), .O(po103));
  buf  g571(.a(pi015), .O(po104));
  buf  g572(.a(pi064), .O(po105));
  buf  g573(.a(pi009), .O(po106));
  buf  g574(.a(pi102), .O(po107));
  buf  g575(.a(pi011), .O(po108));
  buf  g576(.a(pi007), .O(po109));
  buf  g577(.a(pi013), .O(po110));
endmodule


